
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std .ALL;


entity Comunicator is
Generic(
    -- the ammount of bit to recive
    RECIVING_SIZE: integer := 6144;

    -- the ammount of bit to recive
    SENDING_SIZE: integer := 2048;

    -- the numer of clock cicle the macine wait before sending the data back
    CLOCK_REPLYING_TIMER: integer := 5

);
Port(
    CLK: in std_logic;
    TX: out std_logic;
    RX: in std_logic;
    reset: in std_logic;
    waiting_indicator: out std_logic;
    loading_indicator: out std_logic;
    weating_sending_indicator: out std_logic
);
end Comunicator;

architecture Behavioral of Comunicator is

    Type StateType is (Waiting,Loading,Weating_sending,Weating_sending2,Weating_sending3);

    signal state: StateType := Waiting;

    signal TX_reciver: std_logic := '1';
    signal RX_reciver: std_logic := '1';

    signal TX_transmeater: std_logic := '1';
    signal RX_transmeater: std_logic := '1';


    signal data_ready_reciver:  std_logic := '0';

    signal data_in: std_logic_vector(RECIVING_SIZE-1 downto 0);
    signal data_out: std_logic_vector(SENDING_SIZE-1 downto 0);

    signal transmeater_trigger: std_logic := '0';
    signal transmeater_finishd: std_logic := '0';

    signal counter: unsigned(31 downto 0);

    signal reset_signal:  std_logic := '1';

    signal second_reset:  std_logic := '1';

    -- inputs
    signal input_X0_Y0_r: unsigned(7 downto 0);
signal input_X0_Y0_g: unsigned(7 downto 0);
signal input_X0_Y0_b: unsigned(7 downto 0);
signal input_X0_Y1_r: unsigned(7 downto 0);
signal input_X0_Y1_g: unsigned(7 downto 0);
signal input_X0_Y1_b: unsigned(7 downto 0);
signal input_X0_Y2_r: unsigned(7 downto 0);
signal input_X0_Y2_g: unsigned(7 downto 0);
signal input_X0_Y2_b: unsigned(7 downto 0);
signal input_X0_Y3_r: unsigned(7 downto 0);
signal input_X0_Y3_g: unsigned(7 downto 0);
signal input_X0_Y3_b: unsigned(7 downto 0);
signal input_X0_Y4_r: unsigned(7 downto 0);
signal input_X0_Y4_g: unsigned(7 downto 0);
signal input_X0_Y4_b: unsigned(7 downto 0);
signal input_X0_Y5_r: unsigned(7 downto 0);
signal input_X0_Y5_g: unsigned(7 downto 0);
signal input_X0_Y5_b: unsigned(7 downto 0);
signal input_X0_Y6_r: unsigned(7 downto 0);
signal input_X0_Y6_g: unsigned(7 downto 0);
signal input_X0_Y6_b: unsigned(7 downto 0);
signal input_X0_Y7_r: unsigned(7 downto 0);
signal input_X0_Y7_g: unsigned(7 downto 0);
signal input_X0_Y7_b: unsigned(7 downto 0);
signal input_X0_Y8_r: unsigned(7 downto 0);
signal input_X0_Y8_g: unsigned(7 downto 0);
signal input_X0_Y8_b: unsigned(7 downto 0);
signal input_X0_Y9_r: unsigned(7 downto 0);
signal input_X0_Y9_g: unsigned(7 downto 0);
signal input_X0_Y9_b: unsigned(7 downto 0);
signal input_X0_Y10_r: unsigned(7 downto 0);
signal input_X0_Y10_g: unsigned(7 downto 0);
signal input_X0_Y10_b: unsigned(7 downto 0);
signal input_X0_Y11_r: unsigned(7 downto 0);
signal input_X0_Y11_g: unsigned(7 downto 0);
signal input_X0_Y11_b: unsigned(7 downto 0);
signal input_X0_Y12_r: unsigned(7 downto 0);
signal input_X0_Y12_g: unsigned(7 downto 0);
signal input_X0_Y12_b: unsigned(7 downto 0);
signal input_X0_Y13_r: unsigned(7 downto 0);
signal input_X0_Y13_g: unsigned(7 downto 0);
signal input_X0_Y13_b: unsigned(7 downto 0);
signal input_X0_Y14_r: unsigned(7 downto 0);
signal input_X0_Y14_g: unsigned(7 downto 0);
signal input_X0_Y14_b: unsigned(7 downto 0);
signal input_X0_Y15_r: unsigned(7 downto 0);
signal input_X0_Y15_g: unsigned(7 downto 0);
signal input_X0_Y15_b: unsigned(7 downto 0);
signal input_X1_Y0_r: unsigned(7 downto 0);
signal input_X1_Y0_g: unsigned(7 downto 0);
signal input_X1_Y0_b: unsigned(7 downto 0);
signal input_X1_Y1_r: unsigned(7 downto 0);
signal input_X1_Y1_g: unsigned(7 downto 0);
signal input_X1_Y1_b: unsigned(7 downto 0);
signal input_X1_Y2_r: unsigned(7 downto 0);
signal input_X1_Y2_g: unsigned(7 downto 0);
signal input_X1_Y2_b: unsigned(7 downto 0);
signal input_X1_Y3_r: unsigned(7 downto 0);
signal input_X1_Y3_g: unsigned(7 downto 0);
signal input_X1_Y3_b: unsigned(7 downto 0);
signal input_X1_Y4_r: unsigned(7 downto 0);
signal input_X1_Y4_g: unsigned(7 downto 0);
signal input_X1_Y4_b: unsigned(7 downto 0);
signal input_X1_Y5_r: unsigned(7 downto 0);
signal input_X1_Y5_g: unsigned(7 downto 0);
signal input_X1_Y5_b: unsigned(7 downto 0);
signal input_X1_Y6_r: unsigned(7 downto 0);
signal input_X1_Y6_g: unsigned(7 downto 0);
signal input_X1_Y6_b: unsigned(7 downto 0);
signal input_X1_Y7_r: unsigned(7 downto 0);
signal input_X1_Y7_g: unsigned(7 downto 0);
signal input_X1_Y7_b: unsigned(7 downto 0);
signal input_X1_Y8_r: unsigned(7 downto 0);
signal input_X1_Y8_g: unsigned(7 downto 0);
signal input_X1_Y8_b: unsigned(7 downto 0);
signal input_X1_Y9_r: unsigned(7 downto 0);
signal input_X1_Y9_g: unsigned(7 downto 0);
signal input_X1_Y9_b: unsigned(7 downto 0);
signal input_X1_Y10_r: unsigned(7 downto 0);
signal input_X1_Y10_g: unsigned(7 downto 0);
signal input_X1_Y10_b: unsigned(7 downto 0);
signal input_X1_Y11_r: unsigned(7 downto 0);
signal input_X1_Y11_g: unsigned(7 downto 0);
signal input_X1_Y11_b: unsigned(7 downto 0);
signal input_X1_Y12_r: unsigned(7 downto 0);
signal input_X1_Y12_g: unsigned(7 downto 0);
signal input_X1_Y12_b: unsigned(7 downto 0);
signal input_X1_Y13_r: unsigned(7 downto 0);
signal input_X1_Y13_g: unsigned(7 downto 0);
signal input_X1_Y13_b: unsigned(7 downto 0);
signal input_X1_Y14_r: unsigned(7 downto 0);
signal input_X1_Y14_g: unsigned(7 downto 0);
signal input_X1_Y14_b: unsigned(7 downto 0);
signal input_X1_Y15_r: unsigned(7 downto 0);
signal input_X1_Y15_g: unsigned(7 downto 0);
signal input_X1_Y15_b: unsigned(7 downto 0);
signal input_X2_Y0_r: unsigned(7 downto 0);
signal input_X2_Y0_g: unsigned(7 downto 0);
signal input_X2_Y0_b: unsigned(7 downto 0);
signal input_X2_Y1_r: unsigned(7 downto 0);
signal input_X2_Y1_g: unsigned(7 downto 0);
signal input_X2_Y1_b: unsigned(7 downto 0);
signal input_X2_Y2_r: unsigned(7 downto 0);
signal input_X2_Y2_g: unsigned(7 downto 0);
signal input_X2_Y2_b: unsigned(7 downto 0);
signal input_X2_Y3_r: unsigned(7 downto 0);
signal input_X2_Y3_g: unsigned(7 downto 0);
signal input_X2_Y3_b: unsigned(7 downto 0);
signal input_X2_Y4_r: unsigned(7 downto 0);
signal input_X2_Y4_g: unsigned(7 downto 0);
signal input_X2_Y4_b: unsigned(7 downto 0);
signal input_X2_Y5_r: unsigned(7 downto 0);
signal input_X2_Y5_g: unsigned(7 downto 0);
signal input_X2_Y5_b: unsigned(7 downto 0);
signal input_X2_Y6_r: unsigned(7 downto 0);
signal input_X2_Y6_g: unsigned(7 downto 0);
signal input_X2_Y6_b: unsigned(7 downto 0);
signal input_X2_Y7_r: unsigned(7 downto 0);
signal input_X2_Y7_g: unsigned(7 downto 0);
signal input_X2_Y7_b: unsigned(7 downto 0);
signal input_X2_Y8_r: unsigned(7 downto 0);
signal input_X2_Y8_g: unsigned(7 downto 0);
signal input_X2_Y8_b: unsigned(7 downto 0);
signal input_X2_Y9_r: unsigned(7 downto 0);
signal input_X2_Y9_g: unsigned(7 downto 0);
signal input_X2_Y9_b: unsigned(7 downto 0);
signal input_X2_Y10_r: unsigned(7 downto 0);
signal input_X2_Y10_g: unsigned(7 downto 0);
signal input_X2_Y10_b: unsigned(7 downto 0);
signal input_X2_Y11_r: unsigned(7 downto 0);
signal input_X2_Y11_g: unsigned(7 downto 0);
signal input_X2_Y11_b: unsigned(7 downto 0);
signal input_X2_Y12_r: unsigned(7 downto 0);
signal input_X2_Y12_g: unsigned(7 downto 0);
signal input_X2_Y12_b: unsigned(7 downto 0);
signal input_X2_Y13_r: unsigned(7 downto 0);
signal input_X2_Y13_g: unsigned(7 downto 0);
signal input_X2_Y13_b: unsigned(7 downto 0);
signal input_X2_Y14_r: unsigned(7 downto 0);
signal input_X2_Y14_g: unsigned(7 downto 0);
signal input_X2_Y14_b: unsigned(7 downto 0);
signal input_X2_Y15_r: unsigned(7 downto 0);
signal input_X2_Y15_g: unsigned(7 downto 0);
signal input_X2_Y15_b: unsigned(7 downto 0);
signal input_X3_Y0_r: unsigned(7 downto 0);
signal input_X3_Y0_g: unsigned(7 downto 0);
signal input_X3_Y0_b: unsigned(7 downto 0);
signal input_X3_Y1_r: unsigned(7 downto 0);
signal input_X3_Y1_g: unsigned(7 downto 0);
signal input_X3_Y1_b: unsigned(7 downto 0);
signal input_X3_Y2_r: unsigned(7 downto 0);
signal input_X3_Y2_g: unsigned(7 downto 0);
signal input_X3_Y2_b: unsigned(7 downto 0);
signal input_X3_Y3_r: unsigned(7 downto 0);
signal input_X3_Y3_g: unsigned(7 downto 0);
signal input_X3_Y3_b: unsigned(7 downto 0);
signal input_X3_Y4_r: unsigned(7 downto 0);
signal input_X3_Y4_g: unsigned(7 downto 0);
signal input_X3_Y4_b: unsigned(7 downto 0);
signal input_X3_Y5_r: unsigned(7 downto 0);
signal input_X3_Y5_g: unsigned(7 downto 0);
signal input_X3_Y5_b: unsigned(7 downto 0);
signal input_X3_Y6_r: unsigned(7 downto 0);
signal input_X3_Y6_g: unsigned(7 downto 0);
signal input_X3_Y6_b: unsigned(7 downto 0);
signal input_X3_Y7_r: unsigned(7 downto 0);
signal input_X3_Y7_g: unsigned(7 downto 0);
signal input_X3_Y7_b: unsigned(7 downto 0);
signal input_X3_Y8_r: unsigned(7 downto 0);
signal input_X3_Y8_g: unsigned(7 downto 0);
signal input_X3_Y8_b: unsigned(7 downto 0);
signal input_X3_Y9_r: unsigned(7 downto 0);
signal input_X3_Y9_g: unsigned(7 downto 0);
signal input_X3_Y9_b: unsigned(7 downto 0);
signal input_X3_Y10_r: unsigned(7 downto 0);
signal input_X3_Y10_g: unsigned(7 downto 0);
signal input_X3_Y10_b: unsigned(7 downto 0);
signal input_X3_Y11_r: unsigned(7 downto 0);
signal input_X3_Y11_g: unsigned(7 downto 0);
signal input_X3_Y11_b: unsigned(7 downto 0);
signal input_X3_Y12_r: unsigned(7 downto 0);
signal input_X3_Y12_g: unsigned(7 downto 0);
signal input_X3_Y12_b: unsigned(7 downto 0);
signal input_X3_Y13_r: unsigned(7 downto 0);
signal input_X3_Y13_g: unsigned(7 downto 0);
signal input_X3_Y13_b: unsigned(7 downto 0);
signal input_X3_Y14_r: unsigned(7 downto 0);
signal input_X3_Y14_g: unsigned(7 downto 0);
signal input_X3_Y14_b: unsigned(7 downto 0);
signal input_X3_Y15_r: unsigned(7 downto 0);
signal input_X3_Y15_g: unsigned(7 downto 0);
signal input_X3_Y15_b: unsigned(7 downto 0);
signal input_X4_Y0_r: unsigned(7 downto 0);
signal input_X4_Y0_g: unsigned(7 downto 0);
signal input_X4_Y0_b: unsigned(7 downto 0);
signal input_X4_Y1_r: unsigned(7 downto 0);
signal input_X4_Y1_g: unsigned(7 downto 0);
signal input_X4_Y1_b: unsigned(7 downto 0);
signal input_X4_Y2_r: unsigned(7 downto 0);
signal input_X4_Y2_g: unsigned(7 downto 0);
signal input_X4_Y2_b: unsigned(7 downto 0);
signal input_X4_Y3_r: unsigned(7 downto 0);
signal input_X4_Y3_g: unsigned(7 downto 0);
signal input_X4_Y3_b: unsigned(7 downto 0);
signal input_X4_Y4_r: unsigned(7 downto 0);
signal input_X4_Y4_g: unsigned(7 downto 0);
signal input_X4_Y4_b: unsigned(7 downto 0);
signal input_X4_Y5_r: unsigned(7 downto 0);
signal input_X4_Y5_g: unsigned(7 downto 0);
signal input_X4_Y5_b: unsigned(7 downto 0);
signal input_X4_Y6_r: unsigned(7 downto 0);
signal input_X4_Y6_g: unsigned(7 downto 0);
signal input_X4_Y6_b: unsigned(7 downto 0);
signal input_X4_Y7_r: unsigned(7 downto 0);
signal input_X4_Y7_g: unsigned(7 downto 0);
signal input_X4_Y7_b: unsigned(7 downto 0);
signal input_X4_Y8_r: unsigned(7 downto 0);
signal input_X4_Y8_g: unsigned(7 downto 0);
signal input_X4_Y8_b: unsigned(7 downto 0);
signal input_X4_Y9_r: unsigned(7 downto 0);
signal input_X4_Y9_g: unsigned(7 downto 0);
signal input_X4_Y9_b: unsigned(7 downto 0);
signal input_X4_Y10_r: unsigned(7 downto 0);
signal input_X4_Y10_g: unsigned(7 downto 0);
signal input_X4_Y10_b: unsigned(7 downto 0);
signal input_X4_Y11_r: unsigned(7 downto 0);
signal input_X4_Y11_g: unsigned(7 downto 0);
signal input_X4_Y11_b: unsigned(7 downto 0);
signal input_X4_Y12_r: unsigned(7 downto 0);
signal input_X4_Y12_g: unsigned(7 downto 0);
signal input_X4_Y12_b: unsigned(7 downto 0);
signal input_X4_Y13_r: unsigned(7 downto 0);
signal input_X4_Y13_g: unsigned(7 downto 0);
signal input_X4_Y13_b: unsigned(7 downto 0);
signal input_X4_Y14_r: unsigned(7 downto 0);
signal input_X4_Y14_g: unsigned(7 downto 0);
signal input_X4_Y14_b: unsigned(7 downto 0);
signal input_X4_Y15_r: unsigned(7 downto 0);
signal input_X4_Y15_g: unsigned(7 downto 0);
signal input_X4_Y15_b: unsigned(7 downto 0);
signal input_X5_Y0_r: unsigned(7 downto 0);
signal input_X5_Y0_g: unsigned(7 downto 0);
signal input_X5_Y0_b: unsigned(7 downto 0);
signal input_X5_Y1_r: unsigned(7 downto 0);
signal input_X5_Y1_g: unsigned(7 downto 0);
signal input_X5_Y1_b: unsigned(7 downto 0);
signal input_X5_Y2_r: unsigned(7 downto 0);
signal input_X5_Y2_g: unsigned(7 downto 0);
signal input_X5_Y2_b: unsigned(7 downto 0);
signal input_X5_Y3_r: unsigned(7 downto 0);
signal input_X5_Y3_g: unsigned(7 downto 0);
signal input_X5_Y3_b: unsigned(7 downto 0);
signal input_X5_Y4_r: unsigned(7 downto 0);
signal input_X5_Y4_g: unsigned(7 downto 0);
signal input_X5_Y4_b: unsigned(7 downto 0);
signal input_X5_Y5_r: unsigned(7 downto 0);
signal input_X5_Y5_g: unsigned(7 downto 0);
signal input_X5_Y5_b: unsigned(7 downto 0);
signal input_X5_Y6_r: unsigned(7 downto 0);
signal input_X5_Y6_g: unsigned(7 downto 0);
signal input_X5_Y6_b: unsigned(7 downto 0);
signal input_X5_Y7_r: unsigned(7 downto 0);
signal input_X5_Y7_g: unsigned(7 downto 0);
signal input_X5_Y7_b: unsigned(7 downto 0);
signal input_X5_Y8_r: unsigned(7 downto 0);
signal input_X5_Y8_g: unsigned(7 downto 0);
signal input_X5_Y8_b: unsigned(7 downto 0);
signal input_X5_Y9_r: unsigned(7 downto 0);
signal input_X5_Y9_g: unsigned(7 downto 0);
signal input_X5_Y9_b: unsigned(7 downto 0);
signal input_X5_Y10_r: unsigned(7 downto 0);
signal input_X5_Y10_g: unsigned(7 downto 0);
signal input_X5_Y10_b: unsigned(7 downto 0);
signal input_X5_Y11_r: unsigned(7 downto 0);
signal input_X5_Y11_g: unsigned(7 downto 0);
signal input_X5_Y11_b: unsigned(7 downto 0);
signal input_X5_Y12_r: unsigned(7 downto 0);
signal input_X5_Y12_g: unsigned(7 downto 0);
signal input_X5_Y12_b: unsigned(7 downto 0);
signal input_X5_Y13_r: unsigned(7 downto 0);
signal input_X5_Y13_g: unsigned(7 downto 0);
signal input_X5_Y13_b: unsigned(7 downto 0);
signal input_X5_Y14_r: unsigned(7 downto 0);
signal input_X5_Y14_g: unsigned(7 downto 0);
signal input_X5_Y14_b: unsigned(7 downto 0);
signal input_X5_Y15_r: unsigned(7 downto 0);
signal input_X5_Y15_g: unsigned(7 downto 0);
signal input_X5_Y15_b: unsigned(7 downto 0);
signal input_X6_Y0_r: unsigned(7 downto 0);
signal input_X6_Y0_g: unsigned(7 downto 0);
signal input_X6_Y0_b: unsigned(7 downto 0);
signal input_X6_Y1_r: unsigned(7 downto 0);
signal input_X6_Y1_g: unsigned(7 downto 0);
signal input_X6_Y1_b: unsigned(7 downto 0);
signal input_X6_Y2_r: unsigned(7 downto 0);
signal input_X6_Y2_g: unsigned(7 downto 0);
signal input_X6_Y2_b: unsigned(7 downto 0);
signal input_X6_Y3_r: unsigned(7 downto 0);
signal input_X6_Y3_g: unsigned(7 downto 0);
signal input_X6_Y3_b: unsigned(7 downto 0);
signal input_X6_Y4_r: unsigned(7 downto 0);
signal input_X6_Y4_g: unsigned(7 downto 0);
signal input_X6_Y4_b: unsigned(7 downto 0);
signal input_X6_Y5_r: unsigned(7 downto 0);
signal input_X6_Y5_g: unsigned(7 downto 0);
signal input_X6_Y5_b: unsigned(7 downto 0);
signal input_X6_Y6_r: unsigned(7 downto 0);
signal input_X6_Y6_g: unsigned(7 downto 0);
signal input_X6_Y6_b: unsigned(7 downto 0);
signal input_X6_Y7_r: unsigned(7 downto 0);
signal input_X6_Y7_g: unsigned(7 downto 0);
signal input_X6_Y7_b: unsigned(7 downto 0);
signal input_X6_Y8_r: unsigned(7 downto 0);
signal input_X6_Y8_g: unsigned(7 downto 0);
signal input_X6_Y8_b: unsigned(7 downto 0);
signal input_X6_Y9_r: unsigned(7 downto 0);
signal input_X6_Y9_g: unsigned(7 downto 0);
signal input_X6_Y9_b: unsigned(7 downto 0);
signal input_X6_Y10_r: unsigned(7 downto 0);
signal input_X6_Y10_g: unsigned(7 downto 0);
signal input_X6_Y10_b: unsigned(7 downto 0);
signal input_X6_Y11_r: unsigned(7 downto 0);
signal input_X6_Y11_g: unsigned(7 downto 0);
signal input_X6_Y11_b: unsigned(7 downto 0);
signal input_X6_Y12_r: unsigned(7 downto 0);
signal input_X6_Y12_g: unsigned(7 downto 0);
signal input_X6_Y12_b: unsigned(7 downto 0);
signal input_X6_Y13_r: unsigned(7 downto 0);
signal input_X6_Y13_g: unsigned(7 downto 0);
signal input_X6_Y13_b: unsigned(7 downto 0);
signal input_X6_Y14_r: unsigned(7 downto 0);
signal input_X6_Y14_g: unsigned(7 downto 0);
signal input_X6_Y14_b: unsigned(7 downto 0);
signal input_X6_Y15_r: unsigned(7 downto 0);
signal input_X6_Y15_g: unsigned(7 downto 0);
signal input_X6_Y15_b: unsigned(7 downto 0);
signal input_X7_Y0_r: unsigned(7 downto 0);
signal input_X7_Y0_g: unsigned(7 downto 0);
signal input_X7_Y0_b: unsigned(7 downto 0);
signal input_X7_Y1_r: unsigned(7 downto 0);
signal input_X7_Y1_g: unsigned(7 downto 0);
signal input_X7_Y1_b: unsigned(7 downto 0);
signal input_X7_Y2_r: unsigned(7 downto 0);
signal input_X7_Y2_g: unsigned(7 downto 0);
signal input_X7_Y2_b: unsigned(7 downto 0);
signal input_X7_Y3_r: unsigned(7 downto 0);
signal input_X7_Y3_g: unsigned(7 downto 0);
signal input_X7_Y3_b: unsigned(7 downto 0);
signal input_X7_Y4_r: unsigned(7 downto 0);
signal input_X7_Y4_g: unsigned(7 downto 0);
signal input_X7_Y4_b: unsigned(7 downto 0);
signal input_X7_Y5_r: unsigned(7 downto 0);
signal input_X7_Y5_g: unsigned(7 downto 0);
signal input_X7_Y5_b: unsigned(7 downto 0);
signal input_X7_Y6_r: unsigned(7 downto 0);
signal input_X7_Y6_g: unsigned(7 downto 0);
signal input_X7_Y6_b: unsigned(7 downto 0);
signal input_X7_Y7_r: unsigned(7 downto 0);
signal input_X7_Y7_g: unsigned(7 downto 0);
signal input_X7_Y7_b: unsigned(7 downto 0);
signal input_X7_Y8_r: unsigned(7 downto 0);
signal input_X7_Y8_g: unsigned(7 downto 0);
signal input_X7_Y8_b: unsigned(7 downto 0);
signal input_X7_Y9_r: unsigned(7 downto 0);
signal input_X7_Y9_g: unsigned(7 downto 0);
signal input_X7_Y9_b: unsigned(7 downto 0);
signal input_X7_Y10_r: unsigned(7 downto 0);
signal input_X7_Y10_g: unsigned(7 downto 0);
signal input_X7_Y10_b: unsigned(7 downto 0);
signal input_X7_Y11_r: unsigned(7 downto 0);
signal input_X7_Y11_g: unsigned(7 downto 0);
signal input_X7_Y11_b: unsigned(7 downto 0);
signal input_X7_Y12_r: unsigned(7 downto 0);
signal input_X7_Y12_g: unsigned(7 downto 0);
signal input_X7_Y12_b: unsigned(7 downto 0);
signal input_X7_Y13_r: unsigned(7 downto 0);
signal input_X7_Y13_g: unsigned(7 downto 0);
signal input_X7_Y13_b: unsigned(7 downto 0);
signal input_X7_Y14_r: unsigned(7 downto 0);
signal input_X7_Y14_g: unsigned(7 downto 0);
signal input_X7_Y14_b: unsigned(7 downto 0);
signal input_X7_Y15_r: unsigned(7 downto 0);
signal input_X7_Y15_g: unsigned(7 downto 0);
signal input_X7_Y15_b: unsigned(7 downto 0);
signal input_X8_Y0_r: unsigned(7 downto 0);
signal input_X8_Y0_g: unsigned(7 downto 0);
signal input_X8_Y0_b: unsigned(7 downto 0);
signal input_X8_Y1_r: unsigned(7 downto 0);
signal input_X8_Y1_g: unsigned(7 downto 0);
signal input_X8_Y1_b: unsigned(7 downto 0);
signal input_X8_Y2_r: unsigned(7 downto 0);
signal input_X8_Y2_g: unsigned(7 downto 0);
signal input_X8_Y2_b: unsigned(7 downto 0);
signal input_X8_Y3_r: unsigned(7 downto 0);
signal input_X8_Y3_g: unsigned(7 downto 0);
signal input_X8_Y3_b: unsigned(7 downto 0);
signal input_X8_Y4_r: unsigned(7 downto 0);
signal input_X8_Y4_g: unsigned(7 downto 0);
signal input_X8_Y4_b: unsigned(7 downto 0);
signal input_X8_Y5_r: unsigned(7 downto 0);
signal input_X8_Y5_g: unsigned(7 downto 0);
signal input_X8_Y5_b: unsigned(7 downto 0);
signal input_X8_Y6_r: unsigned(7 downto 0);
signal input_X8_Y6_g: unsigned(7 downto 0);
signal input_X8_Y6_b: unsigned(7 downto 0);
signal input_X8_Y7_r: unsigned(7 downto 0);
signal input_X8_Y7_g: unsigned(7 downto 0);
signal input_X8_Y7_b: unsigned(7 downto 0);
signal input_X8_Y8_r: unsigned(7 downto 0);
signal input_X8_Y8_g: unsigned(7 downto 0);
signal input_X8_Y8_b: unsigned(7 downto 0);
signal input_X8_Y9_r: unsigned(7 downto 0);
signal input_X8_Y9_g: unsigned(7 downto 0);
signal input_X8_Y9_b: unsigned(7 downto 0);
signal input_X8_Y10_r: unsigned(7 downto 0);
signal input_X8_Y10_g: unsigned(7 downto 0);
signal input_X8_Y10_b: unsigned(7 downto 0);
signal input_X8_Y11_r: unsigned(7 downto 0);
signal input_X8_Y11_g: unsigned(7 downto 0);
signal input_X8_Y11_b: unsigned(7 downto 0);
signal input_X8_Y12_r: unsigned(7 downto 0);
signal input_X8_Y12_g: unsigned(7 downto 0);
signal input_X8_Y12_b: unsigned(7 downto 0);
signal input_X8_Y13_r: unsigned(7 downto 0);
signal input_X8_Y13_g: unsigned(7 downto 0);
signal input_X8_Y13_b: unsigned(7 downto 0);
signal input_X8_Y14_r: unsigned(7 downto 0);
signal input_X8_Y14_g: unsigned(7 downto 0);
signal input_X8_Y14_b: unsigned(7 downto 0);
signal input_X8_Y15_r: unsigned(7 downto 0);
signal input_X8_Y15_g: unsigned(7 downto 0);
signal input_X8_Y15_b: unsigned(7 downto 0);
signal input_X9_Y0_r: unsigned(7 downto 0);
signal input_X9_Y0_g: unsigned(7 downto 0);
signal input_X9_Y0_b: unsigned(7 downto 0);
signal input_X9_Y1_r: unsigned(7 downto 0);
signal input_X9_Y1_g: unsigned(7 downto 0);
signal input_X9_Y1_b: unsigned(7 downto 0);
signal input_X9_Y2_r: unsigned(7 downto 0);
signal input_X9_Y2_g: unsigned(7 downto 0);
signal input_X9_Y2_b: unsigned(7 downto 0);
signal input_X9_Y3_r: unsigned(7 downto 0);
signal input_X9_Y3_g: unsigned(7 downto 0);
signal input_X9_Y3_b: unsigned(7 downto 0);
signal input_X9_Y4_r: unsigned(7 downto 0);
signal input_X9_Y4_g: unsigned(7 downto 0);
signal input_X9_Y4_b: unsigned(7 downto 0);
signal input_X9_Y5_r: unsigned(7 downto 0);
signal input_X9_Y5_g: unsigned(7 downto 0);
signal input_X9_Y5_b: unsigned(7 downto 0);
signal input_X9_Y6_r: unsigned(7 downto 0);
signal input_X9_Y6_g: unsigned(7 downto 0);
signal input_X9_Y6_b: unsigned(7 downto 0);
signal input_X9_Y7_r: unsigned(7 downto 0);
signal input_X9_Y7_g: unsigned(7 downto 0);
signal input_X9_Y7_b: unsigned(7 downto 0);
signal input_X9_Y8_r: unsigned(7 downto 0);
signal input_X9_Y8_g: unsigned(7 downto 0);
signal input_X9_Y8_b: unsigned(7 downto 0);
signal input_X9_Y9_r: unsigned(7 downto 0);
signal input_X9_Y9_g: unsigned(7 downto 0);
signal input_X9_Y9_b: unsigned(7 downto 0);
signal input_X9_Y10_r: unsigned(7 downto 0);
signal input_X9_Y10_g: unsigned(7 downto 0);
signal input_X9_Y10_b: unsigned(7 downto 0);
signal input_X9_Y11_r: unsigned(7 downto 0);
signal input_X9_Y11_g: unsigned(7 downto 0);
signal input_X9_Y11_b: unsigned(7 downto 0);
signal input_X9_Y12_r: unsigned(7 downto 0);
signal input_X9_Y12_g: unsigned(7 downto 0);
signal input_X9_Y12_b: unsigned(7 downto 0);
signal input_X9_Y13_r: unsigned(7 downto 0);
signal input_X9_Y13_g: unsigned(7 downto 0);
signal input_X9_Y13_b: unsigned(7 downto 0);
signal input_X9_Y14_r: unsigned(7 downto 0);
signal input_X9_Y14_g: unsigned(7 downto 0);
signal input_X9_Y14_b: unsigned(7 downto 0);
signal input_X9_Y15_r: unsigned(7 downto 0);
signal input_X9_Y15_g: unsigned(7 downto 0);
signal input_X9_Y15_b: unsigned(7 downto 0);
signal input_X10_Y0_r: unsigned(7 downto 0);
signal input_X10_Y0_g: unsigned(7 downto 0);
signal input_X10_Y0_b: unsigned(7 downto 0);
signal input_X10_Y1_r: unsigned(7 downto 0);
signal input_X10_Y1_g: unsigned(7 downto 0);
signal input_X10_Y1_b: unsigned(7 downto 0);
signal input_X10_Y2_r: unsigned(7 downto 0);
signal input_X10_Y2_g: unsigned(7 downto 0);
signal input_X10_Y2_b: unsigned(7 downto 0);
signal input_X10_Y3_r: unsigned(7 downto 0);
signal input_X10_Y3_g: unsigned(7 downto 0);
signal input_X10_Y3_b: unsigned(7 downto 0);
signal input_X10_Y4_r: unsigned(7 downto 0);
signal input_X10_Y4_g: unsigned(7 downto 0);
signal input_X10_Y4_b: unsigned(7 downto 0);
signal input_X10_Y5_r: unsigned(7 downto 0);
signal input_X10_Y5_g: unsigned(7 downto 0);
signal input_X10_Y5_b: unsigned(7 downto 0);
signal input_X10_Y6_r: unsigned(7 downto 0);
signal input_X10_Y6_g: unsigned(7 downto 0);
signal input_X10_Y6_b: unsigned(7 downto 0);
signal input_X10_Y7_r: unsigned(7 downto 0);
signal input_X10_Y7_g: unsigned(7 downto 0);
signal input_X10_Y7_b: unsigned(7 downto 0);
signal input_X10_Y8_r: unsigned(7 downto 0);
signal input_X10_Y8_g: unsigned(7 downto 0);
signal input_X10_Y8_b: unsigned(7 downto 0);
signal input_X10_Y9_r: unsigned(7 downto 0);
signal input_X10_Y9_g: unsigned(7 downto 0);
signal input_X10_Y9_b: unsigned(7 downto 0);
signal input_X10_Y10_r: unsigned(7 downto 0);
signal input_X10_Y10_g: unsigned(7 downto 0);
signal input_X10_Y10_b: unsigned(7 downto 0);
signal input_X10_Y11_r: unsigned(7 downto 0);
signal input_X10_Y11_g: unsigned(7 downto 0);
signal input_X10_Y11_b: unsigned(7 downto 0);
signal input_X10_Y12_r: unsigned(7 downto 0);
signal input_X10_Y12_g: unsigned(7 downto 0);
signal input_X10_Y12_b: unsigned(7 downto 0);
signal input_X10_Y13_r: unsigned(7 downto 0);
signal input_X10_Y13_g: unsigned(7 downto 0);
signal input_X10_Y13_b: unsigned(7 downto 0);
signal input_X10_Y14_r: unsigned(7 downto 0);
signal input_X10_Y14_g: unsigned(7 downto 0);
signal input_X10_Y14_b: unsigned(7 downto 0);
signal input_X10_Y15_r: unsigned(7 downto 0);
signal input_X10_Y15_g: unsigned(7 downto 0);
signal input_X10_Y15_b: unsigned(7 downto 0);
signal input_X11_Y0_r: unsigned(7 downto 0);
signal input_X11_Y0_g: unsigned(7 downto 0);
signal input_X11_Y0_b: unsigned(7 downto 0);
signal input_X11_Y1_r: unsigned(7 downto 0);
signal input_X11_Y1_g: unsigned(7 downto 0);
signal input_X11_Y1_b: unsigned(7 downto 0);
signal input_X11_Y2_r: unsigned(7 downto 0);
signal input_X11_Y2_g: unsigned(7 downto 0);
signal input_X11_Y2_b: unsigned(7 downto 0);
signal input_X11_Y3_r: unsigned(7 downto 0);
signal input_X11_Y3_g: unsigned(7 downto 0);
signal input_X11_Y3_b: unsigned(7 downto 0);
signal input_X11_Y4_r: unsigned(7 downto 0);
signal input_X11_Y4_g: unsigned(7 downto 0);
signal input_X11_Y4_b: unsigned(7 downto 0);
signal input_X11_Y5_r: unsigned(7 downto 0);
signal input_X11_Y5_g: unsigned(7 downto 0);
signal input_X11_Y5_b: unsigned(7 downto 0);
signal input_X11_Y6_r: unsigned(7 downto 0);
signal input_X11_Y6_g: unsigned(7 downto 0);
signal input_X11_Y6_b: unsigned(7 downto 0);
signal input_X11_Y7_r: unsigned(7 downto 0);
signal input_X11_Y7_g: unsigned(7 downto 0);
signal input_X11_Y7_b: unsigned(7 downto 0);
signal input_X11_Y8_r: unsigned(7 downto 0);
signal input_X11_Y8_g: unsigned(7 downto 0);
signal input_X11_Y8_b: unsigned(7 downto 0);
signal input_X11_Y9_r: unsigned(7 downto 0);
signal input_X11_Y9_g: unsigned(7 downto 0);
signal input_X11_Y9_b: unsigned(7 downto 0);
signal input_X11_Y10_r: unsigned(7 downto 0);
signal input_X11_Y10_g: unsigned(7 downto 0);
signal input_X11_Y10_b: unsigned(7 downto 0);
signal input_X11_Y11_r: unsigned(7 downto 0);
signal input_X11_Y11_g: unsigned(7 downto 0);
signal input_X11_Y11_b: unsigned(7 downto 0);
signal input_X11_Y12_r: unsigned(7 downto 0);
signal input_X11_Y12_g: unsigned(7 downto 0);
signal input_X11_Y12_b: unsigned(7 downto 0);
signal input_X11_Y13_r: unsigned(7 downto 0);
signal input_X11_Y13_g: unsigned(7 downto 0);
signal input_X11_Y13_b: unsigned(7 downto 0);
signal input_X11_Y14_r: unsigned(7 downto 0);
signal input_X11_Y14_g: unsigned(7 downto 0);
signal input_X11_Y14_b: unsigned(7 downto 0);
signal input_X11_Y15_r: unsigned(7 downto 0);
signal input_X11_Y15_g: unsigned(7 downto 0);
signal input_X11_Y15_b: unsigned(7 downto 0);
signal input_X12_Y0_r: unsigned(7 downto 0);
signal input_X12_Y0_g: unsigned(7 downto 0);
signal input_X12_Y0_b: unsigned(7 downto 0);
signal input_X12_Y1_r: unsigned(7 downto 0);
signal input_X12_Y1_g: unsigned(7 downto 0);
signal input_X12_Y1_b: unsigned(7 downto 0);
signal input_X12_Y2_r: unsigned(7 downto 0);
signal input_X12_Y2_g: unsigned(7 downto 0);
signal input_X12_Y2_b: unsigned(7 downto 0);
signal input_X12_Y3_r: unsigned(7 downto 0);
signal input_X12_Y3_g: unsigned(7 downto 0);
signal input_X12_Y3_b: unsigned(7 downto 0);
signal input_X12_Y4_r: unsigned(7 downto 0);
signal input_X12_Y4_g: unsigned(7 downto 0);
signal input_X12_Y4_b: unsigned(7 downto 0);
signal input_X12_Y5_r: unsigned(7 downto 0);
signal input_X12_Y5_g: unsigned(7 downto 0);
signal input_X12_Y5_b: unsigned(7 downto 0);
signal input_X12_Y6_r: unsigned(7 downto 0);
signal input_X12_Y6_g: unsigned(7 downto 0);
signal input_X12_Y6_b: unsigned(7 downto 0);
signal input_X12_Y7_r: unsigned(7 downto 0);
signal input_X12_Y7_g: unsigned(7 downto 0);
signal input_X12_Y7_b: unsigned(7 downto 0);
signal input_X12_Y8_r: unsigned(7 downto 0);
signal input_X12_Y8_g: unsigned(7 downto 0);
signal input_X12_Y8_b: unsigned(7 downto 0);
signal input_X12_Y9_r: unsigned(7 downto 0);
signal input_X12_Y9_g: unsigned(7 downto 0);
signal input_X12_Y9_b: unsigned(7 downto 0);
signal input_X12_Y10_r: unsigned(7 downto 0);
signal input_X12_Y10_g: unsigned(7 downto 0);
signal input_X12_Y10_b: unsigned(7 downto 0);
signal input_X12_Y11_r: unsigned(7 downto 0);
signal input_X12_Y11_g: unsigned(7 downto 0);
signal input_X12_Y11_b: unsigned(7 downto 0);
signal input_X12_Y12_r: unsigned(7 downto 0);
signal input_X12_Y12_g: unsigned(7 downto 0);
signal input_X12_Y12_b: unsigned(7 downto 0);
signal input_X12_Y13_r: unsigned(7 downto 0);
signal input_X12_Y13_g: unsigned(7 downto 0);
signal input_X12_Y13_b: unsigned(7 downto 0);
signal input_X12_Y14_r: unsigned(7 downto 0);
signal input_X12_Y14_g: unsigned(7 downto 0);
signal input_X12_Y14_b: unsigned(7 downto 0);
signal input_X12_Y15_r: unsigned(7 downto 0);
signal input_X12_Y15_g: unsigned(7 downto 0);
signal input_X12_Y15_b: unsigned(7 downto 0);
signal input_X13_Y0_r: unsigned(7 downto 0);
signal input_X13_Y0_g: unsigned(7 downto 0);
signal input_X13_Y0_b: unsigned(7 downto 0);
signal input_X13_Y1_r: unsigned(7 downto 0);
signal input_X13_Y1_g: unsigned(7 downto 0);
signal input_X13_Y1_b: unsigned(7 downto 0);
signal input_X13_Y2_r: unsigned(7 downto 0);
signal input_X13_Y2_g: unsigned(7 downto 0);
signal input_X13_Y2_b: unsigned(7 downto 0);
signal input_X13_Y3_r: unsigned(7 downto 0);
signal input_X13_Y3_g: unsigned(7 downto 0);
signal input_X13_Y3_b: unsigned(7 downto 0);
signal input_X13_Y4_r: unsigned(7 downto 0);
signal input_X13_Y4_g: unsigned(7 downto 0);
signal input_X13_Y4_b: unsigned(7 downto 0);
signal input_X13_Y5_r: unsigned(7 downto 0);
signal input_X13_Y5_g: unsigned(7 downto 0);
signal input_X13_Y5_b: unsigned(7 downto 0);
signal input_X13_Y6_r: unsigned(7 downto 0);
signal input_X13_Y6_g: unsigned(7 downto 0);
signal input_X13_Y6_b: unsigned(7 downto 0);
signal input_X13_Y7_r: unsigned(7 downto 0);
signal input_X13_Y7_g: unsigned(7 downto 0);
signal input_X13_Y7_b: unsigned(7 downto 0);
signal input_X13_Y8_r: unsigned(7 downto 0);
signal input_X13_Y8_g: unsigned(7 downto 0);
signal input_X13_Y8_b: unsigned(7 downto 0);
signal input_X13_Y9_r: unsigned(7 downto 0);
signal input_X13_Y9_g: unsigned(7 downto 0);
signal input_X13_Y9_b: unsigned(7 downto 0);
signal input_X13_Y10_r: unsigned(7 downto 0);
signal input_X13_Y10_g: unsigned(7 downto 0);
signal input_X13_Y10_b: unsigned(7 downto 0);
signal input_X13_Y11_r: unsigned(7 downto 0);
signal input_X13_Y11_g: unsigned(7 downto 0);
signal input_X13_Y11_b: unsigned(7 downto 0);
signal input_X13_Y12_r: unsigned(7 downto 0);
signal input_X13_Y12_g: unsigned(7 downto 0);
signal input_X13_Y12_b: unsigned(7 downto 0);
signal input_X13_Y13_r: unsigned(7 downto 0);
signal input_X13_Y13_g: unsigned(7 downto 0);
signal input_X13_Y13_b: unsigned(7 downto 0);
signal input_X13_Y14_r: unsigned(7 downto 0);
signal input_X13_Y14_g: unsigned(7 downto 0);
signal input_X13_Y14_b: unsigned(7 downto 0);
signal input_X13_Y15_r: unsigned(7 downto 0);
signal input_X13_Y15_g: unsigned(7 downto 0);
signal input_X13_Y15_b: unsigned(7 downto 0);
signal input_X14_Y0_r: unsigned(7 downto 0);
signal input_X14_Y0_g: unsigned(7 downto 0);
signal input_X14_Y0_b: unsigned(7 downto 0);
signal input_X14_Y1_r: unsigned(7 downto 0);
signal input_X14_Y1_g: unsigned(7 downto 0);
signal input_X14_Y1_b: unsigned(7 downto 0);
signal input_X14_Y2_r: unsigned(7 downto 0);
signal input_X14_Y2_g: unsigned(7 downto 0);
signal input_X14_Y2_b: unsigned(7 downto 0);
signal input_X14_Y3_r: unsigned(7 downto 0);
signal input_X14_Y3_g: unsigned(7 downto 0);
signal input_X14_Y3_b: unsigned(7 downto 0);
signal input_X14_Y4_r: unsigned(7 downto 0);
signal input_X14_Y4_g: unsigned(7 downto 0);
signal input_X14_Y4_b: unsigned(7 downto 0);
signal input_X14_Y5_r: unsigned(7 downto 0);
signal input_X14_Y5_g: unsigned(7 downto 0);
signal input_X14_Y5_b: unsigned(7 downto 0);
signal input_X14_Y6_r: unsigned(7 downto 0);
signal input_X14_Y6_g: unsigned(7 downto 0);
signal input_X14_Y6_b: unsigned(7 downto 0);
signal input_X14_Y7_r: unsigned(7 downto 0);
signal input_X14_Y7_g: unsigned(7 downto 0);
signal input_X14_Y7_b: unsigned(7 downto 0);
signal input_X14_Y8_r: unsigned(7 downto 0);
signal input_X14_Y8_g: unsigned(7 downto 0);
signal input_X14_Y8_b: unsigned(7 downto 0);
signal input_X14_Y9_r: unsigned(7 downto 0);
signal input_X14_Y9_g: unsigned(7 downto 0);
signal input_X14_Y9_b: unsigned(7 downto 0);
signal input_X14_Y10_r: unsigned(7 downto 0);
signal input_X14_Y10_g: unsigned(7 downto 0);
signal input_X14_Y10_b: unsigned(7 downto 0);
signal input_X14_Y11_r: unsigned(7 downto 0);
signal input_X14_Y11_g: unsigned(7 downto 0);
signal input_X14_Y11_b: unsigned(7 downto 0);
signal input_X14_Y12_r: unsigned(7 downto 0);
signal input_X14_Y12_g: unsigned(7 downto 0);
signal input_X14_Y12_b: unsigned(7 downto 0);
signal input_X14_Y13_r: unsigned(7 downto 0);
signal input_X14_Y13_g: unsigned(7 downto 0);
signal input_X14_Y13_b: unsigned(7 downto 0);
signal input_X14_Y14_r: unsigned(7 downto 0);
signal input_X14_Y14_g: unsigned(7 downto 0);
signal input_X14_Y14_b: unsigned(7 downto 0);
signal input_X14_Y15_r: unsigned(7 downto 0);
signal input_X14_Y15_g: unsigned(7 downto 0);
signal input_X14_Y15_b: unsigned(7 downto 0);
signal input_X15_Y0_r: unsigned(7 downto 0);
signal input_X15_Y0_g: unsigned(7 downto 0);
signal input_X15_Y0_b: unsigned(7 downto 0);
signal input_X15_Y1_r: unsigned(7 downto 0);
signal input_X15_Y1_g: unsigned(7 downto 0);
signal input_X15_Y1_b: unsigned(7 downto 0);
signal input_X15_Y2_r: unsigned(7 downto 0);
signal input_X15_Y2_g: unsigned(7 downto 0);
signal input_X15_Y2_b: unsigned(7 downto 0);
signal input_X15_Y3_r: unsigned(7 downto 0);
signal input_X15_Y3_g: unsigned(7 downto 0);
signal input_X15_Y3_b: unsigned(7 downto 0);
signal input_X15_Y4_r: unsigned(7 downto 0);
signal input_X15_Y4_g: unsigned(7 downto 0);
signal input_X15_Y4_b: unsigned(7 downto 0);
signal input_X15_Y5_r: unsigned(7 downto 0);
signal input_X15_Y5_g: unsigned(7 downto 0);
signal input_X15_Y5_b: unsigned(7 downto 0);
signal input_X15_Y6_r: unsigned(7 downto 0);
signal input_X15_Y6_g: unsigned(7 downto 0);
signal input_X15_Y6_b: unsigned(7 downto 0);
signal input_X15_Y7_r: unsigned(7 downto 0);
signal input_X15_Y7_g: unsigned(7 downto 0);
signal input_X15_Y7_b: unsigned(7 downto 0);
signal input_X15_Y8_r: unsigned(7 downto 0);
signal input_X15_Y8_g: unsigned(7 downto 0);
signal input_X15_Y8_b: unsigned(7 downto 0);
signal input_X15_Y9_r: unsigned(7 downto 0);
signal input_X15_Y9_g: unsigned(7 downto 0);
signal input_X15_Y9_b: unsigned(7 downto 0);
signal input_X15_Y10_r: unsigned(7 downto 0);
signal input_X15_Y10_g: unsigned(7 downto 0);
signal input_X15_Y10_b: unsigned(7 downto 0);
signal input_X15_Y11_r: unsigned(7 downto 0);
signal input_X15_Y11_g: unsigned(7 downto 0);
signal input_X15_Y11_b: unsigned(7 downto 0);
signal input_X15_Y12_r: unsigned(7 downto 0);
signal input_X15_Y12_g: unsigned(7 downto 0);
signal input_X15_Y12_b: unsigned(7 downto 0);
signal input_X15_Y13_r: unsigned(7 downto 0);
signal input_X15_Y13_g: unsigned(7 downto 0);
signal input_X15_Y13_b: unsigned(7 downto 0);
signal input_X15_Y14_r: unsigned(7 downto 0);
signal input_X15_Y14_g: unsigned(7 downto 0);
signal input_X15_Y14_b: unsigned(7 downto 0);
signal input_X15_Y15_r: unsigned(7 downto 0);
signal input_X15_Y15_g: unsigned(7 downto 0);
signal input_X15_Y15_b: unsigned(7 downto 0);


    --output
    signal output_X0_Y0_gray: unsigned(7 downto 0);
signal output_X0_Y1_gray: unsigned(7 downto 0);
signal output_X0_Y2_gray: unsigned(7 downto 0);
signal output_X0_Y3_gray: unsigned(7 downto 0);
signal output_X0_Y4_gray: unsigned(7 downto 0);
signal output_X0_Y5_gray: unsigned(7 downto 0);
signal output_X0_Y6_gray: unsigned(7 downto 0);
signal output_X0_Y7_gray: unsigned(7 downto 0);
signal output_X0_Y8_gray: unsigned(7 downto 0);
signal output_X0_Y9_gray: unsigned(7 downto 0);
signal output_X0_Y10_gray: unsigned(7 downto 0);
signal output_X0_Y11_gray: unsigned(7 downto 0);
signal output_X0_Y12_gray: unsigned(7 downto 0);
signal output_X0_Y13_gray: unsigned(7 downto 0);
signal output_X0_Y14_gray: unsigned(7 downto 0);
signal output_X0_Y15_gray: unsigned(7 downto 0);
signal output_X1_Y0_gray: unsigned(7 downto 0);
signal output_X1_Y1_gray: unsigned(7 downto 0);
signal output_X1_Y2_gray: unsigned(7 downto 0);
signal output_X1_Y3_gray: unsigned(7 downto 0);
signal output_X1_Y4_gray: unsigned(7 downto 0);
signal output_X1_Y5_gray: unsigned(7 downto 0);
signal output_X1_Y6_gray: unsigned(7 downto 0);
signal output_X1_Y7_gray: unsigned(7 downto 0);
signal output_X1_Y8_gray: unsigned(7 downto 0);
signal output_X1_Y9_gray: unsigned(7 downto 0);
signal output_X1_Y10_gray: unsigned(7 downto 0);
signal output_X1_Y11_gray: unsigned(7 downto 0);
signal output_X1_Y12_gray: unsigned(7 downto 0);
signal output_X1_Y13_gray: unsigned(7 downto 0);
signal output_X1_Y14_gray: unsigned(7 downto 0);
signal output_X1_Y15_gray: unsigned(7 downto 0);
signal output_X2_Y0_gray: unsigned(7 downto 0);
signal output_X2_Y1_gray: unsigned(7 downto 0);
signal output_X2_Y2_gray: unsigned(7 downto 0);
signal output_X2_Y3_gray: unsigned(7 downto 0);
signal output_X2_Y4_gray: unsigned(7 downto 0);
signal output_X2_Y5_gray: unsigned(7 downto 0);
signal output_X2_Y6_gray: unsigned(7 downto 0);
signal output_X2_Y7_gray: unsigned(7 downto 0);
signal output_X2_Y8_gray: unsigned(7 downto 0);
signal output_X2_Y9_gray: unsigned(7 downto 0);
signal output_X2_Y10_gray: unsigned(7 downto 0);
signal output_X2_Y11_gray: unsigned(7 downto 0);
signal output_X2_Y12_gray: unsigned(7 downto 0);
signal output_X2_Y13_gray: unsigned(7 downto 0);
signal output_X2_Y14_gray: unsigned(7 downto 0);
signal output_X2_Y15_gray: unsigned(7 downto 0);
signal output_X3_Y0_gray: unsigned(7 downto 0);
signal output_X3_Y1_gray: unsigned(7 downto 0);
signal output_X3_Y2_gray: unsigned(7 downto 0);
signal output_X3_Y3_gray: unsigned(7 downto 0);
signal output_X3_Y4_gray: unsigned(7 downto 0);
signal output_X3_Y5_gray: unsigned(7 downto 0);
signal output_X3_Y6_gray: unsigned(7 downto 0);
signal output_X3_Y7_gray: unsigned(7 downto 0);
signal output_X3_Y8_gray: unsigned(7 downto 0);
signal output_X3_Y9_gray: unsigned(7 downto 0);
signal output_X3_Y10_gray: unsigned(7 downto 0);
signal output_X3_Y11_gray: unsigned(7 downto 0);
signal output_X3_Y12_gray: unsigned(7 downto 0);
signal output_X3_Y13_gray: unsigned(7 downto 0);
signal output_X3_Y14_gray: unsigned(7 downto 0);
signal output_X3_Y15_gray: unsigned(7 downto 0);
signal output_X4_Y0_gray: unsigned(7 downto 0);
signal output_X4_Y1_gray: unsigned(7 downto 0);
signal output_X4_Y2_gray: unsigned(7 downto 0);
signal output_X4_Y3_gray: unsigned(7 downto 0);
signal output_X4_Y4_gray: unsigned(7 downto 0);
signal output_X4_Y5_gray: unsigned(7 downto 0);
signal output_X4_Y6_gray: unsigned(7 downto 0);
signal output_X4_Y7_gray: unsigned(7 downto 0);
signal output_X4_Y8_gray: unsigned(7 downto 0);
signal output_X4_Y9_gray: unsigned(7 downto 0);
signal output_X4_Y10_gray: unsigned(7 downto 0);
signal output_X4_Y11_gray: unsigned(7 downto 0);
signal output_X4_Y12_gray: unsigned(7 downto 0);
signal output_X4_Y13_gray: unsigned(7 downto 0);
signal output_X4_Y14_gray: unsigned(7 downto 0);
signal output_X4_Y15_gray: unsigned(7 downto 0);
signal output_X5_Y0_gray: unsigned(7 downto 0);
signal output_X5_Y1_gray: unsigned(7 downto 0);
signal output_X5_Y2_gray: unsigned(7 downto 0);
signal output_X5_Y3_gray: unsigned(7 downto 0);
signal output_X5_Y4_gray: unsigned(7 downto 0);
signal output_X5_Y5_gray: unsigned(7 downto 0);
signal output_X5_Y6_gray: unsigned(7 downto 0);
signal output_X5_Y7_gray: unsigned(7 downto 0);
signal output_X5_Y8_gray: unsigned(7 downto 0);
signal output_X5_Y9_gray: unsigned(7 downto 0);
signal output_X5_Y10_gray: unsigned(7 downto 0);
signal output_X5_Y11_gray: unsigned(7 downto 0);
signal output_X5_Y12_gray: unsigned(7 downto 0);
signal output_X5_Y13_gray: unsigned(7 downto 0);
signal output_X5_Y14_gray: unsigned(7 downto 0);
signal output_X5_Y15_gray: unsigned(7 downto 0);
signal output_X6_Y0_gray: unsigned(7 downto 0);
signal output_X6_Y1_gray: unsigned(7 downto 0);
signal output_X6_Y2_gray: unsigned(7 downto 0);
signal output_X6_Y3_gray: unsigned(7 downto 0);
signal output_X6_Y4_gray: unsigned(7 downto 0);
signal output_X6_Y5_gray: unsigned(7 downto 0);
signal output_X6_Y6_gray: unsigned(7 downto 0);
signal output_X6_Y7_gray: unsigned(7 downto 0);
signal output_X6_Y8_gray: unsigned(7 downto 0);
signal output_X6_Y9_gray: unsigned(7 downto 0);
signal output_X6_Y10_gray: unsigned(7 downto 0);
signal output_X6_Y11_gray: unsigned(7 downto 0);
signal output_X6_Y12_gray: unsigned(7 downto 0);
signal output_X6_Y13_gray: unsigned(7 downto 0);
signal output_X6_Y14_gray: unsigned(7 downto 0);
signal output_X6_Y15_gray: unsigned(7 downto 0);
signal output_X7_Y0_gray: unsigned(7 downto 0);
signal output_X7_Y1_gray: unsigned(7 downto 0);
signal output_X7_Y2_gray: unsigned(7 downto 0);
signal output_X7_Y3_gray: unsigned(7 downto 0);
signal output_X7_Y4_gray: unsigned(7 downto 0);
signal output_X7_Y5_gray: unsigned(7 downto 0);
signal output_X7_Y6_gray: unsigned(7 downto 0);
signal output_X7_Y7_gray: unsigned(7 downto 0);
signal output_X7_Y8_gray: unsigned(7 downto 0);
signal output_X7_Y9_gray: unsigned(7 downto 0);
signal output_X7_Y10_gray: unsigned(7 downto 0);
signal output_X7_Y11_gray: unsigned(7 downto 0);
signal output_X7_Y12_gray: unsigned(7 downto 0);
signal output_X7_Y13_gray: unsigned(7 downto 0);
signal output_X7_Y14_gray: unsigned(7 downto 0);
signal output_X7_Y15_gray: unsigned(7 downto 0);
signal output_X8_Y0_gray: unsigned(7 downto 0);
signal output_X8_Y1_gray: unsigned(7 downto 0);
signal output_X8_Y2_gray: unsigned(7 downto 0);
signal output_X8_Y3_gray: unsigned(7 downto 0);
signal output_X8_Y4_gray: unsigned(7 downto 0);
signal output_X8_Y5_gray: unsigned(7 downto 0);
signal output_X8_Y6_gray: unsigned(7 downto 0);
signal output_X8_Y7_gray: unsigned(7 downto 0);
signal output_X8_Y8_gray: unsigned(7 downto 0);
signal output_X8_Y9_gray: unsigned(7 downto 0);
signal output_X8_Y10_gray: unsigned(7 downto 0);
signal output_X8_Y11_gray: unsigned(7 downto 0);
signal output_X8_Y12_gray: unsigned(7 downto 0);
signal output_X8_Y13_gray: unsigned(7 downto 0);
signal output_X8_Y14_gray: unsigned(7 downto 0);
signal output_X8_Y15_gray: unsigned(7 downto 0);
signal output_X9_Y0_gray: unsigned(7 downto 0);
signal output_X9_Y1_gray: unsigned(7 downto 0);
signal output_X9_Y2_gray: unsigned(7 downto 0);
signal output_X9_Y3_gray: unsigned(7 downto 0);
signal output_X9_Y4_gray: unsigned(7 downto 0);
signal output_X9_Y5_gray: unsigned(7 downto 0);
signal output_X9_Y6_gray: unsigned(7 downto 0);
signal output_X9_Y7_gray: unsigned(7 downto 0);
signal output_X9_Y8_gray: unsigned(7 downto 0);
signal output_X9_Y9_gray: unsigned(7 downto 0);
signal output_X9_Y10_gray: unsigned(7 downto 0);
signal output_X9_Y11_gray: unsigned(7 downto 0);
signal output_X9_Y12_gray: unsigned(7 downto 0);
signal output_X9_Y13_gray: unsigned(7 downto 0);
signal output_X9_Y14_gray: unsigned(7 downto 0);
signal output_X9_Y15_gray: unsigned(7 downto 0);
signal output_X10_Y0_gray: unsigned(7 downto 0);
signal output_X10_Y1_gray: unsigned(7 downto 0);
signal output_X10_Y2_gray: unsigned(7 downto 0);
signal output_X10_Y3_gray: unsigned(7 downto 0);
signal output_X10_Y4_gray: unsigned(7 downto 0);
signal output_X10_Y5_gray: unsigned(7 downto 0);
signal output_X10_Y6_gray: unsigned(7 downto 0);
signal output_X10_Y7_gray: unsigned(7 downto 0);
signal output_X10_Y8_gray: unsigned(7 downto 0);
signal output_X10_Y9_gray: unsigned(7 downto 0);
signal output_X10_Y10_gray: unsigned(7 downto 0);
signal output_X10_Y11_gray: unsigned(7 downto 0);
signal output_X10_Y12_gray: unsigned(7 downto 0);
signal output_X10_Y13_gray: unsigned(7 downto 0);
signal output_X10_Y14_gray: unsigned(7 downto 0);
signal output_X10_Y15_gray: unsigned(7 downto 0);
signal output_X11_Y0_gray: unsigned(7 downto 0);
signal output_X11_Y1_gray: unsigned(7 downto 0);
signal output_X11_Y2_gray: unsigned(7 downto 0);
signal output_X11_Y3_gray: unsigned(7 downto 0);
signal output_X11_Y4_gray: unsigned(7 downto 0);
signal output_X11_Y5_gray: unsigned(7 downto 0);
signal output_X11_Y6_gray: unsigned(7 downto 0);
signal output_X11_Y7_gray: unsigned(7 downto 0);
signal output_X11_Y8_gray: unsigned(7 downto 0);
signal output_X11_Y9_gray: unsigned(7 downto 0);
signal output_X11_Y10_gray: unsigned(7 downto 0);
signal output_X11_Y11_gray: unsigned(7 downto 0);
signal output_X11_Y12_gray: unsigned(7 downto 0);
signal output_X11_Y13_gray: unsigned(7 downto 0);
signal output_X11_Y14_gray: unsigned(7 downto 0);
signal output_X11_Y15_gray: unsigned(7 downto 0);
signal output_X12_Y0_gray: unsigned(7 downto 0);
signal output_X12_Y1_gray: unsigned(7 downto 0);
signal output_X12_Y2_gray: unsigned(7 downto 0);
signal output_X12_Y3_gray: unsigned(7 downto 0);
signal output_X12_Y4_gray: unsigned(7 downto 0);
signal output_X12_Y5_gray: unsigned(7 downto 0);
signal output_X12_Y6_gray: unsigned(7 downto 0);
signal output_X12_Y7_gray: unsigned(7 downto 0);
signal output_X12_Y8_gray: unsigned(7 downto 0);
signal output_X12_Y9_gray: unsigned(7 downto 0);
signal output_X12_Y10_gray: unsigned(7 downto 0);
signal output_X12_Y11_gray: unsigned(7 downto 0);
signal output_X12_Y12_gray: unsigned(7 downto 0);
signal output_X12_Y13_gray: unsigned(7 downto 0);
signal output_X12_Y14_gray: unsigned(7 downto 0);
signal output_X12_Y15_gray: unsigned(7 downto 0);
signal output_X13_Y0_gray: unsigned(7 downto 0);
signal output_X13_Y1_gray: unsigned(7 downto 0);
signal output_X13_Y2_gray: unsigned(7 downto 0);
signal output_X13_Y3_gray: unsigned(7 downto 0);
signal output_X13_Y4_gray: unsigned(7 downto 0);
signal output_X13_Y5_gray: unsigned(7 downto 0);
signal output_X13_Y6_gray: unsigned(7 downto 0);
signal output_X13_Y7_gray: unsigned(7 downto 0);
signal output_X13_Y8_gray: unsigned(7 downto 0);
signal output_X13_Y9_gray: unsigned(7 downto 0);
signal output_X13_Y10_gray: unsigned(7 downto 0);
signal output_X13_Y11_gray: unsigned(7 downto 0);
signal output_X13_Y12_gray: unsigned(7 downto 0);
signal output_X13_Y13_gray: unsigned(7 downto 0);
signal output_X13_Y14_gray: unsigned(7 downto 0);
signal output_X13_Y15_gray: unsigned(7 downto 0);
signal output_X14_Y0_gray: unsigned(7 downto 0);
signal output_X14_Y1_gray: unsigned(7 downto 0);
signal output_X14_Y2_gray: unsigned(7 downto 0);
signal output_X14_Y3_gray: unsigned(7 downto 0);
signal output_X14_Y4_gray: unsigned(7 downto 0);
signal output_X14_Y5_gray: unsigned(7 downto 0);
signal output_X14_Y6_gray: unsigned(7 downto 0);
signal output_X14_Y7_gray: unsigned(7 downto 0);
signal output_X14_Y8_gray: unsigned(7 downto 0);
signal output_X14_Y9_gray: unsigned(7 downto 0);
signal output_X14_Y10_gray: unsigned(7 downto 0);
signal output_X14_Y11_gray: unsigned(7 downto 0);
signal output_X14_Y12_gray: unsigned(7 downto 0);
signal output_X14_Y13_gray: unsigned(7 downto 0);
signal output_X14_Y14_gray: unsigned(7 downto 0);
signal output_X14_Y15_gray: unsigned(7 downto 0);
signal output_X15_Y0_gray: unsigned(7 downto 0);
signal output_X15_Y1_gray: unsigned(7 downto 0);
signal output_X15_Y2_gray: unsigned(7 downto 0);
signal output_X15_Y3_gray: unsigned(7 downto 0);
signal output_X15_Y4_gray: unsigned(7 downto 0);
signal output_X15_Y5_gray: unsigned(7 downto 0);
signal output_X15_Y6_gray: unsigned(7 downto 0);
signal output_X15_Y7_gray: unsigned(7 downto 0);
signal output_X15_Y8_gray: unsigned(7 downto 0);
signal output_X15_Y9_gray: unsigned(7 downto 0);
signal output_X15_Y10_gray: unsigned(7 downto 0);
signal output_X15_Y11_gray: unsigned(7 downto 0);
signal output_X15_Y12_gray: unsigned(7 downto 0);
signal output_X15_Y13_gray: unsigned(7 downto 0);
signal output_X15_Y14_gray: unsigned(7 downto 0);
signal output_X15_Y15_gray: unsigned(7 downto 0);


begin

    transmeater: entity work.SafeTransmeater
        Generic map(
            RECIVING_SIZE =>  SENDING_SIZE
        )
        port map(
          CLK => CLK,
          TX =>TX_transmeater,
          RX =>RX_transmeater,
          reset =>reset_signal,
          input_trigger => transmeater_trigger,
          input =>data_out,
          send_finished => transmeater_finishd
        );

    reciver: entity work.SafeReciver
        Generic map(
            RECIVING_SIZE =>  RECIVING_SIZE
        )
        port map(
            CLK => CLK,
            RX => RX_reciver,
            TX => TX_reciver,
            reset => reset_signal,
            output_ready => data_ready_reciver,
            output => data_in
        );


    --TX <= TX_reciver when state = Waiting else TX_transmeater;
    TX <= TX_reciver and TX_transmeater;


    RX_reciver <= RX when state = Waiting else '1';
    RX_transmeater <= '1' when state = Waiting else RX;

    waiting_indicator <= '1' when state = Waiting else '0';
    loading_indicator <= '1' when state = Loading else '0';
    weating_sending_indicator <= '1' when state = Weating_sending else '0';

    reset_signal <= reset and second_reset;

    main: process(CLK,reset) begin


        if reset = '0' then
            state <= Waiting;
        end if;

        if rising_edge(CLK) then

            if state = Waiting then
                second_reset <= '1';
                if data_ready_reciver = '1' then
                    state <= Loading;
                    counter <= TO_UNSIGNED(0,32);
                end if;

            elsif state = Loading then
                counter <= counter+1;

                if counter >  TO_UNSIGNED(CLOCK_REPLYING_TIMER,32)then
                    transmeater_trigger <= '1';
                end if;

                if counter >  TO_UNSIGNED(CLOCK_REPLYING_TIMER+2,32)then
                    transmeater_trigger <= '0';
                end if;

                if counter >  TO_UNSIGNED(CLOCK_REPLYING_TIMER+4,32)then
                    state <= Weating_sending;
                end if;


            elsif state = Weating_sending then
                if transmeater_finishd = '1' then
                    state <= Weating_sending2;
                    second_reset <= '0';
                end if;

            elsif state = Weating_sending2 then
                    state <= Weating_sending3;
            elsif state = Weating_sending3 then
                    state <= Waiting;
            end if;


        end if;

    end process;

    --constructing inputs
    input_X0_Y0_r <= unsigned(data_in(7 downto 0));
input_X0_Y0_g <= unsigned(data_in(15 downto 8));
input_X0_Y0_b <= unsigned(data_in(23 downto 16));
input_X0_Y1_r <= unsigned(data_in(31 downto 24));
input_X0_Y1_g <= unsigned(data_in(39 downto 32));
input_X0_Y1_b <= unsigned(data_in(47 downto 40));
input_X0_Y2_r <= unsigned(data_in(55 downto 48));
input_X0_Y2_g <= unsigned(data_in(63 downto 56));
input_X0_Y2_b <= unsigned(data_in(71 downto 64));
input_X0_Y3_r <= unsigned(data_in(79 downto 72));
input_X0_Y3_g <= unsigned(data_in(87 downto 80));
input_X0_Y3_b <= unsigned(data_in(95 downto 88));
input_X0_Y4_r <= unsigned(data_in(103 downto 96));
input_X0_Y4_g <= unsigned(data_in(111 downto 104));
input_X0_Y4_b <= unsigned(data_in(119 downto 112));
input_X0_Y5_r <= unsigned(data_in(127 downto 120));
input_X0_Y5_g <= unsigned(data_in(135 downto 128));
input_X0_Y5_b <= unsigned(data_in(143 downto 136));
input_X0_Y6_r <= unsigned(data_in(151 downto 144));
input_X0_Y6_g <= unsigned(data_in(159 downto 152));
input_X0_Y6_b <= unsigned(data_in(167 downto 160));
input_X0_Y7_r <= unsigned(data_in(175 downto 168));
input_X0_Y7_g <= unsigned(data_in(183 downto 176));
input_X0_Y7_b <= unsigned(data_in(191 downto 184));
input_X0_Y8_r <= unsigned(data_in(199 downto 192));
input_X0_Y8_g <= unsigned(data_in(207 downto 200));
input_X0_Y8_b <= unsigned(data_in(215 downto 208));
input_X0_Y9_r <= unsigned(data_in(223 downto 216));
input_X0_Y9_g <= unsigned(data_in(231 downto 224));
input_X0_Y9_b <= unsigned(data_in(239 downto 232));
input_X0_Y10_r <= unsigned(data_in(247 downto 240));
input_X0_Y10_g <= unsigned(data_in(255 downto 248));
input_X0_Y10_b <= unsigned(data_in(263 downto 256));
input_X0_Y11_r <= unsigned(data_in(271 downto 264));
input_X0_Y11_g <= unsigned(data_in(279 downto 272));
input_X0_Y11_b <= unsigned(data_in(287 downto 280));
input_X0_Y12_r <= unsigned(data_in(295 downto 288));
input_X0_Y12_g <= unsigned(data_in(303 downto 296));
input_X0_Y12_b <= unsigned(data_in(311 downto 304));
input_X0_Y13_r <= unsigned(data_in(319 downto 312));
input_X0_Y13_g <= unsigned(data_in(327 downto 320));
input_X0_Y13_b <= unsigned(data_in(335 downto 328));
input_X0_Y14_r <= unsigned(data_in(343 downto 336));
input_X0_Y14_g <= unsigned(data_in(351 downto 344));
input_X0_Y14_b <= unsigned(data_in(359 downto 352));
input_X0_Y15_r <= unsigned(data_in(367 downto 360));
input_X0_Y15_g <= unsigned(data_in(375 downto 368));
input_X0_Y15_b <= unsigned(data_in(383 downto 376));
input_X1_Y0_r <= unsigned(data_in(391 downto 384));
input_X1_Y0_g <= unsigned(data_in(399 downto 392));
input_X1_Y0_b <= unsigned(data_in(407 downto 400));
input_X1_Y1_r <= unsigned(data_in(415 downto 408));
input_X1_Y1_g <= unsigned(data_in(423 downto 416));
input_X1_Y1_b <= unsigned(data_in(431 downto 424));
input_X1_Y2_r <= unsigned(data_in(439 downto 432));
input_X1_Y2_g <= unsigned(data_in(447 downto 440));
input_X1_Y2_b <= unsigned(data_in(455 downto 448));
input_X1_Y3_r <= unsigned(data_in(463 downto 456));
input_X1_Y3_g <= unsigned(data_in(471 downto 464));
input_X1_Y3_b <= unsigned(data_in(479 downto 472));
input_X1_Y4_r <= unsigned(data_in(487 downto 480));
input_X1_Y4_g <= unsigned(data_in(495 downto 488));
input_X1_Y4_b <= unsigned(data_in(503 downto 496));
input_X1_Y5_r <= unsigned(data_in(511 downto 504));
input_X1_Y5_g <= unsigned(data_in(519 downto 512));
input_X1_Y5_b <= unsigned(data_in(527 downto 520));
input_X1_Y6_r <= unsigned(data_in(535 downto 528));
input_X1_Y6_g <= unsigned(data_in(543 downto 536));
input_X1_Y6_b <= unsigned(data_in(551 downto 544));
input_X1_Y7_r <= unsigned(data_in(559 downto 552));
input_X1_Y7_g <= unsigned(data_in(567 downto 560));
input_X1_Y7_b <= unsigned(data_in(575 downto 568));
input_X1_Y8_r <= unsigned(data_in(583 downto 576));
input_X1_Y8_g <= unsigned(data_in(591 downto 584));
input_X1_Y8_b <= unsigned(data_in(599 downto 592));
input_X1_Y9_r <= unsigned(data_in(607 downto 600));
input_X1_Y9_g <= unsigned(data_in(615 downto 608));
input_X1_Y9_b <= unsigned(data_in(623 downto 616));
input_X1_Y10_r <= unsigned(data_in(631 downto 624));
input_X1_Y10_g <= unsigned(data_in(639 downto 632));
input_X1_Y10_b <= unsigned(data_in(647 downto 640));
input_X1_Y11_r <= unsigned(data_in(655 downto 648));
input_X1_Y11_g <= unsigned(data_in(663 downto 656));
input_X1_Y11_b <= unsigned(data_in(671 downto 664));
input_X1_Y12_r <= unsigned(data_in(679 downto 672));
input_X1_Y12_g <= unsigned(data_in(687 downto 680));
input_X1_Y12_b <= unsigned(data_in(695 downto 688));
input_X1_Y13_r <= unsigned(data_in(703 downto 696));
input_X1_Y13_g <= unsigned(data_in(711 downto 704));
input_X1_Y13_b <= unsigned(data_in(719 downto 712));
input_X1_Y14_r <= unsigned(data_in(727 downto 720));
input_X1_Y14_g <= unsigned(data_in(735 downto 728));
input_X1_Y14_b <= unsigned(data_in(743 downto 736));
input_X1_Y15_r <= unsigned(data_in(751 downto 744));
input_X1_Y15_g <= unsigned(data_in(759 downto 752));
input_X1_Y15_b <= unsigned(data_in(767 downto 760));
input_X2_Y0_r <= unsigned(data_in(775 downto 768));
input_X2_Y0_g <= unsigned(data_in(783 downto 776));
input_X2_Y0_b <= unsigned(data_in(791 downto 784));
input_X2_Y1_r <= unsigned(data_in(799 downto 792));
input_X2_Y1_g <= unsigned(data_in(807 downto 800));
input_X2_Y1_b <= unsigned(data_in(815 downto 808));
input_X2_Y2_r <= unsigned(data_in(823 downto 816));
input_X2_Y2_g <= unsigned(data_in(831 downto 824));
input_X2_Y2_b <= unsigned(data_in(839 downto 832));
input_X2_Y3_r <= unsigned(data_in(847 downto 840));
input_X2_Y3_g <= unsigned(data_in(855 downto 848));
input_X2_Y3_b <= unsigned(data_in(863 downto 856));
input_X2_Y4_r <= unsigned(data_in(871 downto 864));
input_X2_Y4_g <= unsigned(data_in(879 downto 872));
input_X2_Y4_b <= unsigned(data_in(887 downto 880));
input_X2_Y5_r <= unsigned(data_in(895 downto 888));
input_X2_Y5_g <= unsigned(data_in(903 downto 896));
input_X2_Y5_b <= unsigned(data_in(911 downto 904));
input_X2_Y6_r <= unsigned(data_in(919 downto 912));
input_X2_Y6_g <= unsigned(data_in(927 downto 920));
input_X2_Y6_b <= unsigned(data_in(935 downto 928));
input_X2_Y7_r <= unsigned(data_in(943 downto 936));
input_X2_Y7_g <= unsigned(data_in(951 downto 944));
input_X2_Y7_b <= unsigned(data_in(959 downto 952));
input_X2_Y8_r <= unsigned(data_in(967 downto 960));
input_X2_Y8_g <= unsigned(data_in(975 downto 968));
input_X2_Y8_b <= unsigned(data_in(983 downto 976));
input_X2_Y9_r <= unsigned(data_in(991 downto 984));
input_X2_Y9_g <= unsigned(data_in(999 downto 992));
input_X2_Y9_b <= unsigned(data_in(1007 downto 1000));
input_X2_Y10_r <= unsigned(data_in(1015 downto 1008));
input_X2_Y10_g <= unsigned(data_in(1023 downto 1016));
input_X2_Y10_b <= unsigned(data_in(1031 downto 1024));
input_X2_Y11_r <= unsigned(data_in(1039 downto 1032));
input_X2_Y11_g <= unsigned(data_in(1047 downto 1040));
input_X2_Y11_b <= unsigned(data_in(1055 downto 1048));
input_X2_Y12_r <= unsigned(data_in(1063 downto 1056));
input_X2_Y12_g <= unsigned(data_in(1071 downto 1064));
input_X2_Y12_b <= unsigned(data_in(1079 downto 1072));
input_X2_Y13_r <= unsigned(data_in(1087 downto 1080));
input_X2_Y13_g <= unsigned(data_in(1095 downto 1088));
input_X2_Y13_b <= unsigned(data_in(1103 downto 1096));
input_X2_Y14_r <= unsigned(data_in(1111 downto 1104));
input_X2_Y14_g <= unsigned(data_in(1119 downto 1112));
input_X2_Y14_b <= unsigned(data_in(1127 downto 1120));
input_X2_Y15_r <= unsigned(data_in(1135 downto 1128));
input_X2_Y15_g <= unsigned(data_in(1143 downto 1136));
input_X2_Y15_b <= unsigned(data_in(1151 downto 1144));
input_X3_Y0_r <= unsigned(data_in(1159 downto 1152));
input_X3_Y0_g <= unsigned(data_in(1167 downto 1160));
input_X3_Y0_b <= unsigned(data_in(1175 downto 1168));
input_X3_Y1_r <= unsigned(data_in(1183 downto 1176));
input_X3_Y1_g <= unsigned(data_in(1191 downto 1184));
input_X3_Y1_b <= unsigned(data_in(1199 downto 1192));
input_X3_Y2_r <= unsigned(data_in(1207 downto 1200));
input_X3_Y2_g <= unsigned(data_in(1215 downto 1208));
input_X3_Y2_b <= unsigned(data_in(1223 downto 1216));
input_X3_Y3_r <= unsigned(data_in(1231 downto 1224));
input_X3_Y3_g <= unsigned(data_in(1239 downto 1232));
input_X3_Y3_b <= unsigned(data_in(1247 downto 1240));
input_X3_Y4_r <= unsigned(data_in(1255 downto 1248));
input_X3_Y4_g <= unsigned(data_in(1263 downto 1256));
input_X3_Y4_b <= unsigned(data_in(1271 downto 1264));
input_X3_Y5_r <= unsigned(data_in(1279 downto 1272));
input_X3_Y5_g <= unsigned(data_in(1287 downto 1280));
input_X3_Y5_b <= unsigned(data_in(1295 downto 1288));
input_X3_Y6_r <= unsigned(data_in(1303 downto 1296));
input_X3_Y6_g <= unsigned(data_in(1311 downto 1304));
input_X3_Y6_b <= unsigned(data_in(1319 downto 1312));
input_X3_Y7_r <= unsigned(data_in(1327 downto 1320));
input_X3_Y7_g <= unsigned(data_in(1335 downto 1328));
input_X3_Y7_b <= unsigned(data_in(1343 downto 1336));
input_X3_Y8_r <= unsigned(data_in(1351 downto 1344));
input_X3_Y8_g <= unsigned(data_in(1359 downto 1352));
input_X3_Y8_b <= unsigned(data_in(1367 downto 1360));
input_X3_Y9_r <= unsigned(data_in(1375 downto 1368));
input_X3_Y9_g <= unsigned(data_in(1383 downto 1376));
input_X3_Y9_b <= unsigned(data_in(1391 downto 1384));
input_X3_Y10_r <= unsigned(data_in(1399 downto 1392));
input_X3_Y10_g <= unsigned(data_in(1407 downto 1400));
input_X3_Y10_b <= unsigned(data_in(1415 downto 1408));
input_X3_Y11_r <= unsigned(data_in(1423 downto 1416));
input_X3_Y11_g <= unsigned(data_in(1431 downto 1424));
input_X3_Y11_b <= unsigned(data_in(1439 downto 1432));
input_X3_Y12_r <= unsigned(data_in(1447 downto 1440));
input_X3_Y12_g <= unsigned(data_in(1455 downto 1448));
input_X3_Y12_b <= unsigned(data_in(1463 downto 1456));
input_X3_Y13_r <= unsigned(data_in(1471 downto 1464));
input_X3_Y13_g <= unsigned(data_in(1479 downto 1472));
input_X3_Y13_b <= unsigned(data_in(1487 downto 1480));
input_X3_Y14_r <= unsigned(data_in(1495 downto 1488));
input_X3_Y14_g <= unsigned(data_in(1503 downto 1496));
input_X3_Y14_b <= unsigned(data_in(1511 downto 1504));
input_X3_Y15_r <= unsigned(data_in(1519 downto 1512));
input_X3_Y15_g <= unsigned(data_in(1527 downto 1520));
input_X3_Y15_b <= unsigned(data_in(1535 downto 1528));
input_X4_Y0_r <= unsigned(data_in(1543 downto 1536));
input_X4_Y0_g <= unsigned(data_in(1551 downto 1544));
input_X4_Y0_b <= unsigned(data_in(1559 downto 1552));
input_X4_Y1_r <= unsigned(data_in(1567 downto 1560));
input_X4_Y1_g <= unsigned(data_in(1575 downto 1568));
input_X4_Y1_b <= unsigned(data_in(1583 downto 1576));
input_X4_Y2_r <= unsigned(data_in(1591 downto 1584));
input_X4_Y2_g <= unsigned(data_in(1599 downto 1592));
input_X4_Y2_b <= unsigned(data_in(1607 downto 1600));
input_X4_Y3_r <= unsigned(data_in(1615 downto 1608));
input_X4_Y3_g <= unsigned(data_in(1623 downto 1616));
input_X4_Y3_b <= unsigned(data_in(1631 downto 1624));
input_X4_Y4_r <= unsigned(data_in(1639 downto 1632));
input_X4_Y4_g <= unsigned(data_in(1647 downto 1640));
input_X4_Y4_b <= unsigned(data_in(1655 downto 1648));
input_X4_Y5_r <= unsigned(data_in(1663 downto 1656));
input_X4_Y5_g <= unsigned(data_in(1671 downto 1664));
input_X4_Y5_b <= unsigned(data_in(1679 downto 1672));
input_X4_Y6_r <= unsigned(data_in(1687 downto 1680));
input_X4_Y6_g <= unsigned(data_in(1695 downto 1688));
input_X4_Y6_b <= unsigned(data_in(1703 downto 1696));
input_X4_Y7_r <= unsigned(data_in(1711 downto 1704));
input_X4_Y7_g <= unsigned(data_in(1719 downto 1712));
input_X4_Y7_b <= unsigned(data_in(1727 downto 1720));
input_X4_Y8_r <= unsigned(data_in(1735 downto 1728));
input_X4_Y8_g <= unsigned(data_in(1743 downto 1736));
input_X4_Y8_b <= unsigned(data_in(1751 downto 1744));
input_X4_Y9_r <= unsigned(data_in(1759 downto 1752));
input_X4_Y9_g <= unsigned(data_in(1767 downto 1760));
input_X4_Y9_b <= unsigned(data_in(1775 downto 1768));
input_X4_Y10_r <= unsigned(data_in(1783 downto 1776));
input_X4_Y10_g <= unsigned(data_in(1791 downto 1784));
input_X4_Y10_b <= unsigned(data_in(1799 downto 1792));
input_X4_Y11_r <= unsigned(data_in(1807 downto 1800));
input_X4_Y11_g <= unsigned(data_in(1815 downto 1808));
input_X4_Y11_b <= unsigned(data_in(1823 downto 1816));
input_X4_Y12_r <= unsigned(data_in(1831 downto 1824));
input_X4_Y12_g <= unsigned(data_in(1839 downto 1832));
input_X4_Y12_b <= unsigned(data_in(1847 downto 1840));
input_X4_Y13_r <= unsigned(data_in(1855 downto 1848));
input_X4_Y13_g <= unsigned(data_in(1863 downto 1856));
input_X4_Y13_b <= unsigned(data_in(1871 downto 1864));
input_X4_Y14_r <= unsigned(data_in(1879 downto 1872));
input_X4_Y14_g <= unsigned(data_in(1887 downto 1880));
input_X4_Y14_b <= unsigned(data_in(1895 downto 1888));
input_X4_Y15_r <= unsigned(data_in(1903 downto 1896));
input_X4_Y15_g <= unsigned(data_in(1911 downto 1904));
input_X4_Y15_b <= unsigned(data_in(1919 downto 1912));
input_X5_Y0_r <= unsigned(data_in(1927 downto 1920));
input_X5_Y0_g <= unsigned(data_in(1935 downto 1928));
input_X5_Y0_b <= unsigned(data_in(1943 downto 1936));
input_X5_Y1_r <= unsigned(data_in(1951 downto 1944));
input_X5_Y1_g <= unsigned(data_in(1959 downto 1952));
input_X5_Y1_b <= unsigned(data_in(1967 downto 1960));
input_X5_Y2_r <= unsigned(data_in(1975 downto 1968));
input_X5_Y2_g <= unsigned(data_in(1983 downto 1976));
input_X5_Y2_b <= unsigned(data_in(1991 downto 1984));
input_X5_Y3_r <= unsigned(data_in(1999 downto 1992));
input_X5_Y3_g <= unsigned(data_in(2007 downto 2000));
input_X5_Y3_b <= unsigned(data_in(2015 downto 2008));
input_X5_Y4_r <= unsigned(data_in(2023 downto 2016));
input_X5_Y4_g <= unsigned(data_in(2031 downto 2024));
input_X5_Y4_b <= unsigned(data_in(2039 downto 2032));
input_X5_Y5_r <= unsigned(data_in(2047 downto 2040));
input_X5_Y5_g <= unsigned(data_in(2055 downto 2048));
input_X5_Y5_b <= unsigned(data_in(2063 downto 2056));
input_X5_Y6_r <= unsigned(data_in(2071 downto 2064));
input_X5_Y6_g <= unsigned(data_in(2079 downto 2072));
input_X5_Y6_b <= unsigned(data_in(2087 downto 2080));
input_X5_Y7_r <= unsigned(data_in(2095 downto 2088));
input_X5_Y7_g <= unsigned(data_in(2103 downto 2096));
input_X5_Y7_b <= unsigned(data_in(2111 downto 2104));
input_X5_Y8_r <= unsigned(data_in(2119 downto 2112));
input_X5_Y8_g <= unsigned(data_in(2127 downto 2120));
input_X5_Y8_b <= unsigned(data_in(2135 downto 2128));
input_X5_Y9_r <= unsigned(data_in(2143 downto 2136));
input_X5_Y9_g <= unsigned(data_in(2151 downto 2144));
input_X5_Y9_b <= unsigned(data_in(2159 downto 2152));
input_X5_Y10_r <= unsigned(data_in(2167 downto 2160));
input_X5_Y10_g <= unsigned(data_in(2175 downto 2168));
input_X5_Y10_b <= unsigned(data_in(2183 downto 2176));
input_X5_Y11_r <= unsigned(data_in(2191 downto 2184));
input_X5_Y11_g <= unsigned(data_in(2199 downto 2192));
input_X5_Y11_b <= unsigned(data_in(2207 downto 2200));
input_X5_Y12_r <= unsigned(data_in(2215 downto 2208));
input_X5_Y12_g <= unsigned(data_in(2223 downto 2216));
input_X5_Y12_b <= unsigned(data_in(2231 downto 2224));
input_X5_Y13_r <= unsigned(data_in(2239 downto 2232));
input_X5_Y13_g <= unsigned(data_in(2247 downto 2240));
input_X5_Y13_b <= unsigned(data_in(2255 downto 2248));
input_X5_Y14_r <= unsigned(data_in(2263 downto 2256));
input_X5_Y14_g <= unsigned(data_in(2271 downto 2264));
input_X5_Y14_b <= unsigned(data_in(2279 downto 2272));
input_X5_Y15_r <= unsigned(data_in(2287 downto 2280));
input_X5_Y15_g <= unsigned(data_in(2295 downto 2288));
input_X5_Y15_b <= unsigned(data_in(2303 downto 2296));
input_X6_Y0_r <= unsigned(data_in(2311 downto 2304));
input_X6_Y0_g <= unsigned(data_in(2319 downto 2312));
input_X6_Y0_b <= unsigned(data_in(2327 downto 2320));
input_X6_Y1_r <= unsigned(data_in(2335 downto 2328));
input_X6_Y1_g <= unsigned(data_in(2343 downto 2336));
input_X6_Y1_b <= unsigned(data_in(2351 downto 2344));
input_X6_Y2_r <= unsigned(data_in(2359 downto 2352));
input_X6_Y2_g <= unsigned(data_in(2367 downto 2360));
input_X6_Y2_b <= unsigned(data_in(2375 downto 2368));
input_X6_Y3_r <= unsigned(data_in(2383 downto 2376));
input_X6_Y3_g <= unsigned(data_in(2391 downto 2384));
input_X6_Y3_b <= unsigned(data_in(2399 downto 2392));
input_X6_Y4_r <= unsigned(data_in(2407 downto 2400));
input_X6_Y4_g <= unsigned(data_in(2415 downto 2408));
input_X6_Y4_b <= unsigned(data_in(2423 downto 2416));
input_X6_Y5_r <= unsigned(data_in(2431 downto 2424));
input_X6_Y5_g <= unsigned(data_in(2439 downto 2432));
input_X6_Y5_b <= unsigned(data_in(2447 downto 2440));
input_X6_Y6_r <= unsigned(data_in(2455 downto 2448));
input_X6_Y6_g <= unsigned(data_in(2463 downto 2456));
input_X6_Y6_b <= unsigned(data_in(2471 downto 2464));
input_X6_Y7_r <= unsigned(data_in(2479 downto 2472));
input_X6_Y7_g <= unsigned(data_in(2487 downto 2480));
input_X6_Y7_b <= unsigned(data_in(2495 downto 2488));
input_X6_Y8_r <= unsigned(data_in(2503 downto 2496));
input_X6_Y8_g <= unsigned(data_in(2511 downto 2504));
input_X6_Y8_b <= unsigned(data_in(2519 downto 2512));
input_X6_Y9_r <= unsigned(data_in(2527 downto 2520));
input_X6_Y9_g <= unsigned(data_in(2535 downto 2528));
input_X6_Y9_b <= unsigned(data_in(2543 downto 2536));
input_X6_Y10_r <= unsigned(data_in(2551 downto 2544));
input_X6_Y10_g <= unsigned(data_in(2559 downto 2552));
input_X6_Y10_b <= unsigned(data_in(2567 downto 2560));
input_X6_Y11_r <= unsigned(data_in(2575 downto 2568));
input_X6_Y11_g <= unsigned(data_in(2583 downto 2576));
input_X6_Y11_b <= unsigned(data_in(2591 downto 2584));
input_X6_Y12_r <= unsigned(data_in(2599 downto 2592));
input_X6_Y12_g <= unsigned(data_in(2607 downto 2600));
input_X6_Y12_b <= unsigned(data_in(2615 downto 2608));
input_X6_Y13_r <= unsigned(data_in(2623 downto 2616));
input_X6_Y13_g <= unsigned(data_in(2631 downto 2624));
input_X6_Y13_b <= unsigned(data_in(2639 downto 2632));
input_X6_Y14_r <= unsigned(data_in(2647 downto 2640));
input_X6_Y14_g <= unsigned(data_in(2655 downto 2648));
input_X6_Y14_b <= unsigned(data_in(2663 downto 2656));
input_X6_Y15_r <= unsigned(data_in(2671 downto 2664));
input_X6_Y15_g <= unsigned(data_in(2679 downto 2672));
input_X6_Y15_b <= unsigned(data_in(2687 downto 2680));
input_X7_Y0_r <= unsigned(data_in(2695 downto 2688));
input_X7_Y0_g <= unsigned(data_in(2703 downto 2696));
input_X7_Y0_b <= unsigned(data_in(2711 downto 2704));
input_X7_Y1_r <= unsigned(data_in(2719 downto 2712));
input_X7_Y1_g <= unsigned(data_in(2727 downto 2720));
input_X7_Y1_b <= unsigned(data_in(2735 downto 2728));
input_X7_Y2_r <= unsigned(data_in(2743 downto 2736));
input_X7_Y2_g <= unsigned(data_in(2751 downto 2744));
input_X7_Y2_b <= unsigned(data_in(2759 downto 2752));
input_X7_Y3_r <= unsigned(data_in(2767 downto 2760));
input_X7_Y3_g <= unsigned(data_in(2775 downto 2768));
input_X7_Y3_b <= unsigned(data_in(2783 downto 2776));
input_X7_Y4_r <= unsigned(data_in(2791 downto 2784));
input_X7_Y4_g <= unsigned(data_in(2799 downto 2792));
input_X7_Y4_b <= unsigned(data_in(2807 downto 2800));
input_X7_Y5_r <= unsigned(data_in(2815 downto 2808));
input_X7_Y5_g <= unsigned(data_in(2823 downto 2816));
input_X7_Y5_b <= unsigned(data_in(2831 downto 2824));
input_X7_Y6_r <= unsigned(data_in(2839 downto 2832));
input_X7_Y6_g <= unsigned(data_in(2847 downto 2840));
input_X7_Y6_b <= unsigned(data_in(2855 downto 2848));
input_X7_Y7_r <= unsigned(data_in(2863 downto 2856));
input_X7_Y7_g <= unsigned(data_in(2871 downto 2864));
input_X7_Y7_b <= unsigned(data_in(2879 downto 2872));
input_X7_Y8_r <= unsigned(data_in(2887 downto 2880));
input_X7_Y8_g <= unsigned(data_in(2895 downto 2888));
input_X7_Y8_b <= unsigned(data_in(2903 downto 2896));
input_X7_Y9_r <= unsigned(data_in(2911 downto 2904));
input_X7_Y9_g <= unsigned(data_in(2919 downto 2912));
input_X7_Y9_b <= unsigned(data_in(2927 downto 2920));
input_X7_Y10_r <= unsigned(data_in(2935 downto 2928));
input_X7_Y10_g <= unsigned(data_in(2943 downto 2936));
input_X7_Y10_b <= unsigned(data_in(2951 downto 2944));
input_X7_Y11_r <= unsigned(data_in(2959 downto 2952));
input_X7_Y11_g <= unsigned(data_in(2967 downto 2960));
input_X7_Y11_b <= unsigned(data_in(2975 downto 2968));
input_X7_Y12_r <= unsigned(data_in(2983 downto 2976));
input_X7_Y12_g <= unsigned(data_in(2991 downto 2984));
input_X7_Y12_b <= unsigned(data_in(2999 downto 2992));
input_X7_Y13_r <= unsigned(data_in(3007 downto 3000));
input_X7_Y13_g <= unsigned(data_in(3015 downto 3008));
input_X7_Y13_b <= unsigned(data_in(3023 downto 3016));
input_X7_Y14_r <= unsigned(data_in(3031 downto 3024));
input_X7_Y14_g <= unsigned(data_in(3039 downto 3032));
input_X7_Y14_b <= unsigned(data_in(3047 downto 3040));
input_X7_Y15_r <= unsigned(data_in(3055 downto 3048));
input_X7_Y15_g <= unsigned(data_in(3063 downto 3056));
input_X7_Y15_b <= unsigned(data_in(3071 downto 3064));
input_X8_Y0_r <= unsigned(data_in(3079 downto 3072));
input_X8_Y0_g <= unsigned(data_in(3087 downto 3080));
input_X8_Y0_b <= unsigned(data_in(3095 downto 3088));
input_X8_Y1_r <= unsigned(data_in(3103 downto 3096));
input_X8_Y1_g <= unsigned(data_in(3111 downto 3104));
input_X8_Y1_b <= unsigned(data_in(3119 downto 3112));
input_X8_Y2_r <= unsigned(data_in(3127 downto 3120));
input_X8_Y2_g <= unsigned(data_in(3135 downto 3128));
input_X8_Y2_b <= unsigned(data_in(3143 downto 3136));
input_X8_Y3_r <= unsigned(data_in(3151 downto 3144));
input_X8_Y3_g <= unsigned(data_in(3159 downto 3152));
input_X8_Y3_b <= unsigned(data_in(3167 downto 3160));
input_X8_Y4_r <= unsigned(data_in(3175 downto 3168));
input_X8_Y4_g <= unsigned(data_in(3183 downto 3176));
input_X8_Y4_b <= unsigned(data_in(3191 downto 3184));
input_X8_Y5_r <= unsigned(data_in(3199 downto 3192));
input_X8_Y5_g <= unsigned(data_in(3207 downto 3200));
input_X8_Y5_b <= unsigned(data_in(3215 downto 3208));
input_X8_Y6_r <= unsigned(data_in(3223 downto 3216));
input_X8_Y6_g <= unsigned(data_in(3231 downto 3224));
input_X8_Y6_b <= unsigned(data_in(3239 downto 3232));
input_X8_Y7_r <= unsigned(data_in(3247 downto 3240));
input_X8_Y7_g <= unsigned(data_in(3255 downto 3248));
input_X8_Y7_b <= unsigned(data_in(3263 downto 3256));
input_X8_Y8_r <= unsigned(data_in(3271 downto 3264));
input_X8_Y8_g <= unsigned(data_in(3279 downto 3272));
input_X8_Y8_b <= unsigned(data_in(3287 downto 3280));
input_X8_Y9_r <= unsigned(data_in(3295 downto 3288));
input_X8_Y9_g <= unsigned(data_in(3303 downto 3296));
input_X8_Y9_b <= unsigned(data_in(3311 downto 3304));
input_X8_Y10_r <= unsigned(data_in(3319 downto 3312));
input_X8_Y10_g <= unsigned(data_in(3327 downto 3320));
input_X8_Y10_b <= unsigned(data_in(3335 downto 3328));
input_X8_Y11_r <= unsigned(data_in(3343 downto 3336));
input_X8_Y11_g <= unsigned(data_in(3351 downto 3344));
input_X8_Y11_b <= unsigned(data_in(3359 downto 3352));
input_X8_Y12_r <= unsigned(data_in(3367 downto 3360));
input_X8_Y12_g <= unsigned(data_in(3375 downto 3368));
input_X8_Y12_b <= unsigned(data_in(3383 downto 3376));
input_X8_Y13_r <= unsigned(data_in(3391 downto 3384));
input_X8_Y13_g <= unsigned(data_in(3399 downto 3392));
input_X8_Y13_b <= unsigned(data_in(3407 downto 3400));
input_X8_Y14_r <= unsigned(data_in(3415 downto 3408));
input_X8_Y14_g <= unsigned(data_in(3423 downto 3416));
input_X8_Y14_b <= unsigned(data_in(3431 downto 3424));
input_X8_Y15_r <= unsigned(data_in(3439 downto 3432));
input_X8_Y15_g <= unsigned(data_in(3447 downto 3440));
input_X8_Y15_b <= unsigned(data_in(3455 downto 3448));
input_X9_Y0_r <= unsigned(data_in(3463 downto 3456));
input_X9_Y0_g <= unsigned(data_in(3471 downto 3464));
input_X9_Y0_b <= unsigned(data_in(3479 downto 3472));
input_X9_Y1_r <= unsigned(data_in(3487 downto 3480));
input_X9_Y1_g <= unsigned(data_in(3495 downto 3488));
input_X9_Y1_b <= unsigned(data_in(3503 downto 3496));
input_X9_Y2_r <= unsigned(data_in(3511 downto 3504));
input_X9_Y2_g <= unsigned(data_in(3519 downto 3512));
input_X9_Y2_b <= unsigned(data_in(3527 downto 3520));
input_X9_Y3_r <= unsigned(data_in(3535 downto 3528));
input_X9_Y3_g <= unsigned(data_in(3543 downto 3536));
input_X9_Y3_b <= unsigned(data_in(3551 downto 3544));
input_X9_Y4_r <= unsigned(data_in(3559 downto 3552));
input_X9_Y4_g <= unsigned(data_in(3567 downto 3560));
input_X9_Y4_b <= unsigned(data_in(3575 downto 3568));
input_X9_Y5_r <= unsigned(data_in(3583 downto 3576));
input_X9_Y5_g <= unsigned(data_in(3591 downto 3584));
input_X9_Y5_b <= unsigned(data_in(3599 downto 3592));
input_X9_Y6_r <= unsigned(data_in(3607 downto 3600));
input_X9_Y6_g <= unsigned(data_in(3615 downto 3608));
input_X9_Y6_b <= unsigned(data_in(3623 downto 3616));
input_X9_Y7_r <= unsigned(data_in(3631 downto 3624));
input_X9_Y7_g <= unsigned(data_in(3639 downto 3632));
input_X9_Y7_b <= unsigned(data_in(3647 downto 3640));
input_X9_Y8_r <= unsigned(data_in(3655 downto 3648));
input_X9_Y8_g <= unsigned(data_in(3663 downto 3656));
input_X9_Y8_b <= unsigned(data_in(3671 downto 3664));
input_X9_Y9_r <= unsigned(data_in(3679 downto 3672));
input_X9_Y9_g <= unsigned(data_in(3687 downto 3680));
input_X9_Y9_b <= unsigned(data_in(3695 downto 3688));
input_X9_Y10_r <= unsigned(data_in(3703 downto 3696));
input_X9_Y10_g <= unsigned(data_in(3711 downto 3704));
input_X9_Y10_b <= unsigned(data_in(3719 downto 3712));
input_X9_Y11_r <= unsigned(data_in(3727 downto 3720));
input_X9_Y11_g <= unsigned(data_in(3735 downto 3728));
input_X9_Y11_b <= unsigned(data_in(3743 downto 3736));
input_X9_Y12_r <= unsigned(data_in(3751 downto 3744));
input_X9_Y12_g <= unsigned(data_in(3759 downto 3752));
input_X9_Y12_b <= unsigned(data_in(3767 downto 3760));
input_X9_Y13_r <= unsigned(data_in(3775 downto 3768));
input_X9_Y13_g <= unsigned(data_in(3783 downto 3776));
input_X9_Y13_b <= unsigned(data_in(3791 downto 3784));
input_X9_Y14_r <= unsigned(data_in(3799 downto 3792));
input_X9_Y14_g <= unsigned(data_in(3807 downto 3800));
input_X9_Y14_b <= unsigned(data_in(3815 downto 3808));
input_X9_Y15_r <= unsigned(data_in(3823 downto 3816));
input_X9_Y15_g <= unsigned(data_in(3831 downto 3824));
input_X9_Y15_b <= unsigned(data_in(3839 downto 3832));
input_X10_Y0_r <= unsigned(data_in(3847 downto 3840));
input_X10_Y0_g <= unsigned(data_in(3855 downto 3848));
input_X10_Y0_b <= unsigned(data_in(3863 downto 3856));
input_X10_Y1_r <= unsigned(data_in(3871 downto 3864));
input_X10_Y1_g <= unsigned(data_in(3879 downto 3872));
input_X10_Y1_b <= unsigned(data_in(3887 downto 3880));
input_X10_Y2_r <= unsigned(data_in(3895 downto 3888));
input_X10_Y2_g <= unsigned(data_in(3903 downto 3896));
input_X10_Y2_b <= unsigned(data_in(3911 downto 3904));
input_X10_Y3_r <= unsigned(data_in(3919 downto 3912));
input_X10_Y3_g <= unsigned(data_in(3927 downto 3920));
input_X10_Y3_b <= unsigned(data_in(3935 downto 3928));
input_X10_Y4_r <= unsigned(data_in(3943 downto 3936));
input_X10_Y4_g <= unsigned(data_in(3951 downto 3944));
input_X10_Y4_b <= unsigned(data_in(3959 downto 3952));
input_X10_Y5_r <= unsigned(data_in(3967 downto 3960));
input_X10_Y5_g <= unsigned(data_in(3975 downto 3968));
input_X10_Y5_b <= unsigned(data_in(3983 downto 3976));
input_X10_Y6_r <= unsigned(data_in(3991 downto 3984));
input_X10_Y6_g <= unsigned(data_in(3999 downto 3992));
input_X10_Y6_b <= unsigned(data_in(4007 downto 4000));
input_X10_Y7_r <= unsigned(data_in(4015 downto 4008));
input_X10_Y7_g <= unsigned(data_in(4023 downto 4016));
input_X10_Y7_b <= unsigned(data_in(4031 downto 4024));
input_X10_Y8_r <= unsigned(data_in(4039 downto 4032));
input_X10_Y8_g <= unsigned(data_in(4047 downto 4040));
input_X10_Y8_b <= unsigned(data_in(4055 downto 4048));
input_X10_Y9_r <= unsigned(data_in(4063 downto 4056));
input_X10_Y9_g <= unsigned(data_in(4071 downto 4064));
input_X10_Y9_b <= unsigned(data_in(4079 downto 4072));
input_X10_Y10_r <= unsigned(data_in(4087 downto 4080));
input_X10_Y10_g <= unsigned(data_in(4095 downto 4088));
input_X10_Y10_b <= unsigned(data_in(4103 downto 4096));
input_X10_Y11_r <= unsigned(data_in(4111 downto 4104));
input_X10_Y11_g <= unsigned(data_in(4119 downto 4112));
input_X10_Y11_b <= unsigned(data_in(4127 downto 4120));
input_X10_Y12_r <= unsigned(data_in(4135 downto 4128));
input_X10_Y12_g <= unsigned(data_in(4143 downto 4136));
input_X10_Y12_b <= unsigned(data_in(4151 downto 4144));
input_X10_Y13_r <= unsigned(data_in(4159 downto 4152));
input_X10_Y13_g <= unsigned(data_in(4167 downto 4160));
input_X10_Y13_b <= unsigned(data_in(4175 downto 4168));
input_X10_Y14_r <= unsigned(data_in(4183 downto 4176));
input_X10_Y14_g <= unsigned(data_in(4191 downto 4184));
input_X10_Y14_b <= unsigned(data_in(4199 downto 4192));
input_X10_Y15_r <= unsigned(data_in(4207 downto 4200));
input_X10_Y15_g <= unsigned(data_in(4215 downto 4208));
input_X10_Y15_b <= unsigned(data_in(4223 downto 4216));
input_X11_Y0_r <= unsigned(data_in(4231 downto 4224));
input_X11_Y0_g <= unsigned(data_in(4239 downto 4232));
input_X11_Y0_b <= unsigned(data_in(4247 downto 4240));
input_X11_Y1_r <= unsigned(data_in(4255 downto 4248));
input_X11_Y1_g <= unsigned(data_in(4263 downto 4256));
input_X11_Y1_b <= unsigned(data_in(4271 downto 4264));
input_X11_Y2_r <= unsigned(data_in(4279 downto 4272));
input_X11_Y2_g <= unsigned(data_in(4287 downto 4280));
input_X11_Y2_b <= unsigned(data_in(4295 downto 4288));
input_X11_Y3_r <= unsigned(data_in(4303 downto 4296));
input_X11_Y3_g <= unsigned(data_in(4311 downto 4304));
input_X11_Y3_b <= unsigned(data_in(4319 downto 4312));
input_X11_Y4_r <= unsigned(data_in(4327 downto 4320));
input_X11_Y4_g <= unsigned(data_in(4335 downto 4328));
input_X11_Y4_b <= unsigned(data_in(4343 downto 4336));
input_X11_Y5_r <= unsigned(data_in(4351 downto 4344));
input_X11_Y5_g <= unsigned(data_in(4359 downto 4352));
input_X11_Y5_b <= unsigned(data_in(4367 downto 4360));
input_X11_Y6_r <= unsigned(data_in(4375 downto 4368));
input_X11_Y6_g <= unsigned(data_in(4383 downto 4376));
input_X11_Y6_b <= unsigned(data_in(4391 downto 4384));
input_X11_Y7_r <= unsigned(data_in(4399 downto 4392));
input_X11_Y7_g <= unsigned(data_in(4407 downto 4400));
input_X11_Y7_b <= unsigned(data_in(4415 downto 4408));
input_X11_Y8_r <= unsigned(data_in(4423 downto 4416));
input_X11_Y8_g <= unsigned(data_in(4431 downto 4424));
input_X11_Y8_b <= unsigned(data_in(4439 downto 4432));
input_X11_Y9_r <= unsigned(data_in(4447 downto 4440));
input_X11_Y9_g <= unsigned(data_in(4455 downto 4448));
input_X11_Y9_b <= unsigned(data_in(4463 downto 4456));
input_X11_Y10_r <= unsigned(data_in(4471 downto 4464));
input_X11_Y10_g <= unsigned(data_in(4479 downto 4472));
input_X11_Y10_b <= unsigned(data_in(4487 downto 4480));
input_X11_Y11_r <= unsigned(data_in(4495 downto 4488));
input_X11_Y11_g <= unsigned(data_in(4503 downto 4496));
input_X11_Y11_b <= unsigned(data_in(4511 downto 4504));
input_X11_Y12_r <= unsigned(data_in(4519 downto 4512));
input_X11_Y12_g <= unsigned(data_in(4527 downto 4520));
input_X11_Y12_b <= unsigned(data_in(4535 downto 4528));
input_X11_Y13_r <= unsigned(data_in(4543 downto 4536));
input_X11_Y13_g <= unsigned(data_in(4551 downto 4544));
input_X11_Y13_b <= unsigned(data_in(4559 downto 4552));
input_X11_Y14_r <= unsigned(data_in(4567 downto 4560));
input_X11_Y14_g <= unsigned(data_in(4575 downto 4568));
input_X11_Y14_b <= unsigned(data_in(4583 downto 4576));
input_X11_Y15_r <= unsigned(data_in(4591 downto 4584));
input_X11_Y15_g <= unsigned(data_in(4599 downto 4592));
input_X11_Y15_b <= unsigned(data_in(4607 downto 4600));
input_X12_Y0_r <= unsigned(data_in(4615 downto 4608));
input_X12_Y0_g <= unsigned(data_in(4623 downto 4616));
input_X12_Y0_b <= unsigned(data_in(4631 downto 4624));
input_X12_Y1_r <= unsigned(data_in(4639 downto 4632));
input_X12_Y1_g <= unsigned(data_in(4647 downto 4640));
input_X12_Y1_b <= unsigned(data_in(4655 downto 4648));
input_X12_Y2_r <= unsigned(data_in(4663 downto 4656));
input_X12_Y2_g <= unsigned(data_in(4671 downto 4664));
input_X12_Y2_b <= unsigned(data_in(4679 downto 4672));
input_X12_Y3_r <= unsigned(data_in(4687 downto 4680));
input_X12_Y3_g <= unsigned(data_in(4695 downto 4688));
input_X12_Y3_b <= unsigned(data_in(4703 downto 4696));
input_X12_Y4_r <= unsigned(data_in(4711 downto 4704));
input_X12_Y4_g <= unsigned(data_in(4719 downto 4712));
input_X12_Y4_b <= unsigned(data_in(4727 downto 4720));
input_X12_Y5_r <= unsigned(data_in(4735 downto 4728));
input_X12_Y5_g <= unsigned(data_in(4743 downto 4736));
input_X12_Y5_b <= unsigned(data_in(4751 downto 4744));
input_X12_Y6_r <= unsigned(data_in(4759 downto 4752));
input_X12_Y6_g <= unsigned(data_in(4767 downto 4760));
input_X12_Y6_b <= unsigned(data_in(4775 downto 4768));
input_X12_Y7_r <= unsigned(data_in(4783 downto 4776));
input_X12_Y7_g <= unsigned(data_in(4791 downto 4784));
input_X12_Y7_b <= unsigned(data_in(4799 downto 4792));
input_X12_Y8_r <= unsigned(data_in(4807 downto 4800));
input_X12_Y8_g <= unsigned(data_in(4815 downto 4808));
input_X12_Y8_b <= unsigned(data_in(4823 downto 4816));
input_X12_Y9_r <= unsigned(data_in(4831 downto 4824));
input_X12_Y9_g <= unsigned(data_in(4839 downto 4832));
input_X12_Y9_b <= unsigned(data_in(4847 downto 4840));
input_X12_Y10_r <= unsigned(data_in(4855 downto 4848));
input_X12_Y10_g <= unsigned(data_in(4863 downto 4856));
input_X12_Y10_b <= unsigned(data_in(4871 downto 4864));
input_X12_Y11_r <= unsigned(data_in(4879 downto 4872));
input_X12_Y11_g <= unsigned(data_in(4887 downto 4880));
input_X12_Y11_b <= unsigned(data_in(4895 downto 4888));
input_X12_Y12_r <= unsigned(data_in(4903 downto 4896));
input_X12_Y12_g <= unsigned(data_in(4911 downto 4904));
input_X12_Y12_b <= unsigned(data_in(4919 downto 4912));
input_X12_Y13_r <= unsigned(data_in(4927 downto 4920));
input_X12_Y13_g <= unsigned(data_in(4935 downto 4928));
input_X12_Y13_b <= unsigned(data_in(4943 downto 4936));
input_X12_Y14_r <= unsigned(data_in(4951 downto 4944));
input_X12_Y14_g <= unsigned(data_in(4959 downto 4952));
input_X12_Y14_b <= unsigned(data_in(4967 downto 4960));
input_X12_Y15_r <= unsigned(data_in(4975 downto 4968));
input_X12_Y15_g <= unsigned(data_in(4983 downto 4976));
input_X12_Y15_b <= unsigned(data_in(4991 downto 4984));
input_X13_Y0_r <= unsigned(data_in(4999 downto 4992));
input_X13_Y0_g <= unsigned(data_in(5007 downto 5000));
input_X13_Y0_b <= unsigned(data_in(5015 downto 5008));
input_X13_Y1_r <= unsigned(data_in(5023 downto 5016));
input_X13_Y1_g <= unsigned(data_in(5031 downto 5024));
input_X13_Y1_b <= unsigned(data_in(5039 downto 5032));
input_X13_Y2_r <= unsigned(data_in(5047 downto 5040));
input_X13_Y2_g <= unsigned(data_in(5055 downto 5048));
input_X13_Y2_b <= unsigned(data_in(5063 downto 5056));
input_X13_Y3_r <= unsigned(data_in(5071 downto 5064));
input_X13_Y3_g <= unsigned(data_in(5079 downto 5072));
input_X13_Y3_b <= unsigned(data_in(5087 downto 5080));
input_X13_Y4_r <= unsigned(data_in(5095 downto 5088));
input_X13_Y4_g <= unsigned(data_in(5103 downto 5096));
input_X13_Y4_b <= unsigned(data_in(5111 downto 5104));
input_X13_Y5_r <= unsigned(data_in(5119 downto 5112));
input_X13_Y5_g <= unsigned(data_in(5127 downto 5120));
input_X13_Y5_b <= unsigned(data_in(5135 downto 5128));
input_X13_Y6_r <= unsigned(data_in(5143 downto 5136));
input_X13_Y6_g <= unsigned(data_in(5151 downto 5144));
input_X13_Y6_b <= unsigned(data_in(5159 downto 5152));
input_X13_Y7_r <= unsigned(data_in(5167 downto 5160));
input_X13_Y7_g <= unsigned(data_in(5175 downto 5168));
input_X13_Y7_b <= unsigned(data_in(5183 downto 5176));
input_X13_Y8_r <= unsigned(data_in(5191 downto 5184));
input_X13_Y8_g <= unsigned(data_in(5199 downto 5192));
input_X13_Y8_b <= unsigned(data_in(5207 downto 5200));
input_X13_Y9_r <= unsigned(data_in(5215 downto 5208));
input_X13_Y9_g <= unsigned(data_in(5223 downto 5216));
input_X13_Y9_b <= unsigned(data_in(5231 downto 5224));
input_X13_Y10_r <= unsigned(data_in(5239 downto 5232));
input_X13_Y10_g <= unsigned(data_in(5247 downto 5240));
input_X13_Y10_b <= unsigned(data_in(5255 downto 5248));
input_X13_Y11_r <= unsigned(data_in(5263 downto 5256));
input_X13_Y11_g <= unsigned(data_in(5271 downto 5264));
input_X13_Y11_b <= unsigned(data_in(5279 downto 5272));
input_X13_Y12_r <= unsigned(data_in(5287 downto 5280));
input_X13_Y12_g <= unsigned(data_in(5295 downto 5288));
input_X13_Y12_b <= unsigned(data_in(5303 downto 5296));
input_X13_Y13_r <= unsigned(data_in(5311 downto 5304));
input_X13_Y13_g <= unsigned(data_in(5319 downto 5312));
input_X13_Y13_b <= unsigned(data_in(5327 downto 5320));
input_X13_Y14_r <= unsigned(data_in(5335 downto 5328));
input_X13_Y14_g <= unsigned(data_in(5343 downto 5336));
input_X13_Y14_b <= unsigned(data_in(5351 downto 5344));
input_X13_Y15_r <= unsigned(data_in(5359 downto 5352));
input_X13_Y15_g <= unsigned(data_in(5367 downto 5360));
input_X13_Y15_b <= unsigned(data_in(5375 downto 5368));
input_X14_Y0_r <= unsigned(data_in(5383 downto 5376));
input_X14_Y0_g <= unsigned(data_in(5391 downto 5384));
input_X14_Y0_b <= unsigned(data_in(5399 downto 5392));
input_X14_Y1_r <= unsigned(data_in(5407 downto 5400));
input_X14_Y1_g <= unsigned(data_in(5415 downto 5408));
input_X14_Y1_b <= unsigned(data_in(5423 downto 5416));
input_X14_Y2_r <= unsigned(data_in(5431 downto 5424));
input_X14_Y2_g <= unsigned(data_in(5439 downto 5432));
input_X14_Y2_b <= unsigned(data_in(5447 downto 5440));
input_X14_Y3_r <= unsigned(data_in(5455 downto 5448));
input_X14_Y3_g <= unsigned(data_in(5463 downto 5456));
input_X14_Y3_b <= unsigned(data_in(5471 downto 5464));
input_X14_Y4_r <= unsigned(data_in(5479 downto 5472));
input_X14_Y4_g <= unsigned(data_in(5487 downto 5480));
input_X14_Y4_b <= unsigned(data_in(5495 downto 5488));
input_X14_Y5_r <= unsigned(data_in(5503 downto 5496));
input_X14_Y5_g <= unsigned(data_in(5511 downto 5504));
input_X14_Y5_b <= unsigned(data_in(5519 downto 5512));
input_X14_Y6_r <= unsigned(data_in(5527 downto 5520));
input_X14_Y6_g <= unsigned(data_in(5535 downto 5528));
input_X14_Y6_b <= unsigned(data_in(5543 downto 5536));
input_X14_Y7_r <= unsigned(data_in(5551 downto 5544));
input_X14_Y7_g <= unsigned(data_in(5559 downto 5552));
input_X14_Y7_b <= unsigned(data_in(5567 downto 5560));
input_X14_Y8_r <= unsigned(data_in(5575 downto 5568));
input_X14_Y8_g <= unsigned(data_in(5583 downto 5576));
input_X14_Y8_b <= unsigned(data_in(5591 downto 5584));
input_X14_Y9_r <= unsigned(data_in(5599 downto 5592));
input_X14_Y9_g <= unsigned(data_in(5607 downto 5600));
input_X14_Y9_b <= unsigned(data_in(5615 downto 5608));
input_X14_Y10_r <= unsigned(data_in(5623 downto 5616));
input_X14_Y10_g <= unsigned(data_in(5631 downto 5624));
input_X14_Y10_b <= unsigned(data_in(5639 downto 5632));
input_X14_Y11_r <= unsigned(data_in(5647 downto 5640));
input_X14_Y11_g <= unsigned(data_in(5655 downto 5648));
input_X14_Y11_b <= unsigned(data_in(5663 downto 5656));
input_X14_Y12_r <= unsigned(data_in(5671 downto 5664));
input_X14_Y12_g <= unsigned(data_in(5679 downto 5672));
input_X14_Y12_b <= unsigned(data_in(5687 downto 5680));
input_X14_Y13_r <= unsigned(data_in(5695 downto 5688));
input_X14_Y13_g <= unsigned(data_in(5703 downto 5696));
input_X14_Y13_b <= unsigned(data_in(5711 downto 5704));
input_X14_Y14_r <= unsigned(data_in(5719 downto 5712));
input_X14_Y14_g <= unsigned(data_in(5727 downto 5720));
input_X14_Y14_b <= unsigned(data_in(5735 downto 5728));
input_X14_Y15_r <= unsigned(data_in(5743 downto 5736));
input_X14_Y15_g <= unsigned(data_in(5751 downto 5744));
input_X14_Y15_b <= unsigned(data_in(5759 downto 5752));
input_X15_Y0_r <= unsigned(data_in(5767 downto 5760));
input_X15_Y0_g <= unsigned(data_in(5775 downto 5768));
input_X15_Y0_b <= unsigned(data_in(5783 downto 5776));
input_X15_Y1_r <= unsigned(data_in(5791 downto 5784));
input_X15_Y1_g <= unsigned(data_in(5799 downto 5792));
input_X15_Y1_b <= unsigned(data_in(5807 downto 5800));
input_X15_Y2_r <= unsigned(data_in(5815 downto 5808));
input_X15_Y2_g <= unsigned(data_in(5823 downto 5816));
input_X15_Y2_b <= unsigned(data_in(5831 downto 5824));
input_X15_Y3_r <= unsigned(data_in(5839 downto 5832));
input_X15_Y3_g <= unsigned(data_in(5847 downto 5840));
input_X15_Y3_b <= unsigned(data_in(5855 downto 5848));
input_X15_Y4_r <= unsigned(data_in(5863 downto 5856));
input_X15_Y4_g <= unsigned(data_in(5871 downto 5864));
input_X15_Y4_b <= unsigned(data_in(5879 downto 5872));
input_X15_Y5_r <= unsigned(data_in(5887 downto 5880));
input_X15_Y5_g <= unsigned(data_in(5895 downto 5888));
input_X15_Y5_b <= unsigned(data_in(5903 downto 5896));
input_X15_Y6_r <= unsigned(data_in(5911 downto 5904));
input_X15_Y6_g <= unsigned(data_in(5919 downto 5912));
input_X15_Y6_b <= unsigned(data_in(5927 downto 5920));
input_X15_Y7_r <= unsigned(data_in(5935 downto 5928));
input_X15_Y7_g <= unsigned(data_in(5943 downto 5936));
input_X15_Y7_b <= unsigned(data_in(5951 downto 5944));
input_X15_Y8_r <= unsigned(data_in(5959 downto 5952));
input_X15_Y8_g <= unsigned(data_in(5967 downto 5960));
input_X15_Y8_b <= unsigned(data_in(5975 downto 5968));
input_X15_Y9_r <= unsigned(data_in(5983 downto 5976));
input_X15_Y9_g <= unsigned(data_in(5991 downto 5984));
input_X15_Y9_b <= unsigned(data_in(5999 downto 5992));
input_X15_Y10_r <= unsigned(data_in(6007 downto 6000));
input_X15_Y10_g <= unsigned(data_in(6015 downto 6008));
input_X15_Y10_b <= unsigned(data_in(6023 downto 6016));
input_X15_Y11_r <= unsigned(data_in(6031 downto 6024));
input_X15_Y11_g <= unsigned(data_in(6039 downto 6032));
input_X15_Y11_b <= unsigned(data_in(6047 downto 6040));
input_X15_Y12_r <= unsigned(data_in(6055 downto 6048));
input_X15_Y12_g <= unsigned(data_in(6063 downto 6056));
input_X15_Y12_b <= unsigned(data_in(6071 downto 6064));
input_X15_Y13_r <= unsigned(data_in(6079 downto 6072));
input_X15_Y13_g <= unsigned(data_in(6087 downto 6080));
input_X15_Y13_b <= unsigned(data_in(6095 downto 6088));
input_X15_Y14_r <= unsigned(data_in(6103 downto 6096));
input_X15_Y14_g <= unsigned(data_in(6111 downto 6104));
input_X15_Y14_b <= unsigned(data_in(6119 downto 6112));
input_X15_Y15_r <= unsigned(data_in(6127 downto 6120));
input_X15_Y15_g <= unsigned(data_in(6135 downto 6128));
input_X15_Y15_b <= unsigned(data_in(6143 downto 6136));


    --deconstruction outputs
    data_out(7 downto 0) <= std_logic_vector(output_X0_Y0_gray);
data_out(15 downto 8) <= std_logic_vector(output_X0_Y1_gray);
data_out(23 downto 16) <= std_logic_vector(output_X0_Y2_gray);
data_out(31 downto 24) <= std_logic_vector(output_X0_Y3_gray);
data_out(39 downto 32) <= std_logic_vector(output_X0_Y4_gray);
data_out(47 downto 40) <= std_logic_vector(output_X0_Y5_gray);
data_out(55 downto 48) <= std_logic_vector(output_X0_Y6_gray);
data_out(63 downto 56) <= std_logic_vector(output_X0_Y7_gray);
data_out(71 downto 64) <= std_logic_vector(output_X0_Y8_gray);
data_out(79 downto 72) <= std_logic_vector(output_X0_Y9_gray);
data_out(87 downto 80) <= std_logic_vector(output_X0_Y10_gray);
data_out(95 downto 88) <= std_logic_vector(output_X0_Y11_gray);
data_out(103 downto 96) <= std_logic_vector(output_X0_Y12_gray);
data_out(111 downto 104) <= std_logic_vector(output_X0_Y13_gray);
data_out(119 downto 112) <= std_logic_vector(output_X0_Y14_gray);
data_out(127 downto 120) <= std_logic_vector(output_X0_Y15_gray);
data_out(135 downto 128) <= std_logic_vector(output_X1_Y0_gray);
data_out(143 downto 136) <= std_logic_vector(output_X1_Y1_gray);
data_out(151 downto 144) <= std_logic_vector(output_X1_Y2_gray);
data_out(159 downto 152) <= std_logic_vector(output_X1_Y3_gray);
data_out(167 downto 160) <= std_logic_vector(output_X1_Y4_gray);
data_out(175 downto 168) <= std_logic_vector(output_X1_Y5_gray);
data_out(183 downto 176) <= std_logic_vector(output_X1_Y6_gray);
data_out(191 downto 184) <= std_logic_vector(output_X1_Y7_gray);
data_out(199 downto 192) <= std_logic_vector(output_X1_Y8_gray);
data_out(207 downto 200) <= std_logic_vector(output_X1_Y9_gray);
data_out(215 downto 208) <= std_logic_vector(output_X1_Y10_gray);
data_out(223 downto 216) <= std_logic_vector(output_X1_Y11_gray);
data_out(231 downto 224) <= std_logic_vector(output_X1_Y12_gray);
data_out(239 downto 232) <= std_logic_vector(output_X1_Y13_gray);
data_out(247 downto 240) <= std_logic_vector(output_X1_Y14_gray);
data_out(255 downto 248) <= std_logic_vector(output_X1_Y15_gray);
data_out(263 downto 256) <= std_logic_vector(output_X2_Y0_gray);
data_out(271 downto 264) <= std_logic_vector(output_X2_Y1_gray);
data_out(279 downto 272) <= std_logic_vector(output_X2_Y2_gray);
data_out(287 downto 280) <= std_logic_vector(output_X2_Y3_gray);
data_out(295 downto 288) <= std_logic_vector(output_X2_Y4_gray);
data_out(303 downto 296) <= std_logic_vector(output_X2_Y5_gray);
data_out(311 downto 304) <= std_logic_vector(output_X2_Y6_gray);
data_out(319 downto 312) <= std_logic_vector(output_X2_Y7_gray);
data_out(327 downto 320) <= std_logic_vector(output_X2_Y8_gray);
data_out(335 downto 328) <= std_logic_vector(output_X2_Y9_gray);
data_out(343 downto 336) <= std_logic_vector(output_X2_Y10_gray);
data_out(351 downto 344) <= std_logic_vector(output_X2_Y11_gray);
data_out(359 downto 352) <= std_logic_vector(output_X2_Y12_gray);
data_out(367 downto 360) <= std_logic_vector(output_X2_Y13_gray);
data_out(375 downto 368) <= std_logic_vector(output_X2_Y14_gray);
data_out(383 downto 376) <= std_logic_vector(output_X2_Y15_gray);
data_out(391 downto 384) <= std_logic_vector(output_X3_Y0_gray);
data_out(399 downto 392) <= std_logic_vector(output_X3_Y1_gray);
data_out(407 downto 400) <= std_logic_vector(output_X3_Y2_gray);
data_out(415 downto 408) <= std_logic_vector(output_X3_Y3_gray);
data_out(423 downto 416) <= std_logic_vector(output_X3_Y4_gray);
data_out(431 downto 424) <= std_logic_vector(output_X3_Y5_gray);
data_out(439 downto 432) <= std_logic_vector(output_X3_Y6_gray);
data_out(447 downto 440) <= std_logic_vector(output_X3_Y7_gray);
data_out(455 downto 448) <= std_logic_vector(output_X3_Y8_gray);
data_out(463 downto 456) <= std_logic_vector(output_X3_Y9_gray);
data_out(471 downto 464) <= std_logic_vector(output_X3_Y10_gray);
data_out(479 downto 472) <= std_logic_vector(output_X3_Y11_gray);
data_out(487 downto 480) <= std_logic_vector(output_X3_Y12_gray);
data_out(495 downto 488) <= std_logic_vector(output_X3_Y13_gray);
data_out(503 downto 496) <= std_logic_vector(output_X3_Y14_gray);
data_out(511 downto 504) <= std_logic_vector(output_X3_Y15_gray);
data_out(519 downto 512) <= std_logic_vector(output_X4_Y0_gray);
data_out(527 downto 520) <= std_logic_vector(output_X4_Y1_gray);
data_out(535 downto 528) <= std_logic_vector(output_X4_Y2_gray);
data_out(543 downto 536) <= std_logic_vector(output_X4_Y3_gray);
data_out(551 downto 544) <= std_logic_vector(output_X4_Y4_gray);
data_out(559 downto 552) <= std_logic_vector(output_X4_Y5_gray);
data_out(567 downto 560) <= std_logic_vector(output_X4_Y6_gray);
data_out(575 downto 568) <= std_logic_vector(output_X4_Y7_gray);
data_out(583 downto 576) <= std_logic_vector(output_X4_Y8_gray);
data_out(591 downto 584) <= std_logic_vector(output_X4_Y9_gray);
data_out(599 downto 592) <= std_logic_vector(output_X4_Y10_gray);
data_out(607 downto 600) <= std_logic_vector(output_X4_Y11_gray);
data_out(615 downto 608) <= std_logic_vector(output_X4_Y12_gray);
data_out(623 downto 616) <= std_logic_vector(output_X4_Y13_gray);
data_out(631 downto 624) <= std_logic_vector(output_X4_Y14_gray);
data_out(639 downto 632) <= std_logic_vector(output_X4_Y15_gray);
data_out(647 downto 640) <= std_logic_vector(output_X5_Y0_gray);
data_out(655 downto 648) <= std_logic_vector(output_X5_Y1_gray);
data_out(663 downto 656) <= std_logic_vector(output_X5_Y2_gray);
data_out(671 downto 664) <= std_logic_vector(output_X5_Y3_gray);
data_out(679 downto 672) <= std_logic_vector(output_X5_Y4_gray);
data_out(687 downto 680) <= std_logic_vector(output_X5_Y5_gray);
data_out(695 downto 688) <= std_logic_vector(output_X5_Y6_gray);
data_out(703 downto 696) <= std_logic_vector(output_X5_Y7_gray);
data_out(711 downto 704) <= std_logic_vector(output_X5_Y8_gray);
data_out(719 downto 712) <= std_logic_vector(output_X5_Y9_gray);
data_out(727 downto 720) <= std_logic_vector(output_X5_Y10_gray);
data_out(735 downto 728) <= std_logic_vector(output_X5_Y11_gray);
data_out(743 downto 736) <= std_logic_vector(output_X5_Y12_gray);
data_out(751 downto 744) <= std_logic_vector(output_X5_Y13_gray);
data_out(759 downto 752) <= std_logic_vector(output_X5_Y14_gray);
data_out(767 downto 760) <= std_logic_vector(output_X5_Y15_gray);
data_out(775 downto 768) <= std_logic_vector(output_X6_Y0_gray);
data_out(783 downto 776) <= std_logic_vector(output_X6_Y1_gray);
data_out(791 downto 784) <= std_logic_vector(output_X6_Y2_gray);
data_out(799 downto 792) <= std_logic_vector(output_X6_Y3_gray);
data_out(807 downto 800) <= std_logic_vector(output_X6_Y4_gray);
data_out(815 downto 808) <= std_logic_vector(output_X6_Y5_gray);
data_out(823 downto 816) <= std_logic_vector(output_X6_Y6_gray);
data_out(831 downto 824) <= std_logic_vector(output_X6_Y7_gray);
data_out(839 downto 832) <= std_logic_vector(output_X6_Y8_gray);
data_out(847 downto 840) <= std_logic_vector(output_X6_Y9_gray);
data_out(855 downto 848) <= std_logic_vector(output_X6_Y10_gray);
data_out(863 downto 856) <= std_logic_vector(output_X6_Y11_gray);
data_out(871 downto 864) <= std_logic_vector(output_X6_Y12_gray);
data_out(879 downto 872) <= std_logic_vector(output_X6_Y13_gray);
data_out(887 downto 880) <= std_logic_vector(output_X6_Y14_gray);
data_out(895 downto 888) <= std_logic_vector(output_X6_Y15_gray);
data_out(903 downto 896) <= std_logic_vector(output_X7_Y0_gray);
data_out(911 downto 904) <= std_logic_vector(output_X7_Y1_gray);
data_out(919 downto 912) <= std_logic_vector(output_X7_Y2_gray);
data_out(927 downto 920) <= std_logic_vector(output_X7_Y3_gray);
data_out(935 downto 928) <= std_logic_vector(output_X7_Y4_gray);
data_out(943 downto 936) <= std_logic_vector(output_X7_Y5_gray);
data_out(951 downto 944) <= std_logic_vector(output_X7_Y6_gray);
data_out(959 downto 952) <= std_logic_vector(output_X7_Y7_gray);
data_out(967 downto 960) <= std_logic_vector(output_X7_Y8_gray);
data_out(975 downto 968) <= std_logic_vector(output_X7_Y9_gray);
data_out(983 downto 976) <= std_logic_vector(output_X7_Y10_gray);
data_out(991 downto 984) <= std_logic_vector(output_X7_Y11_gray);
data_out(999 downto 992) <= std_logic_vector(output_X7_Y12_gray);
data_out(1007 downto 1000) <= std_logic_vector(output_X7_Y13_gray);
data_out(1015 downto 1008) <= std_logic_vector(output_X7_Y14_gray);
data_out(1023 downto 1016) <= std_logic_vector(output_X7_Y15_gray);
data_out(1031 downto 1024) <= std_logic_vector(output_X8_Y0_gray);
data_out(1039 downto 1032) <= std_logic_vector(output_X8_Y1_gray);
data_out(1047 downto 1040) <= std_logic_vector(output_X8_Y2_gray);
data_out(1055 downto 1048) <= std_logic_vector(output_X8_Y3_gray);
data_out(1063 downto 1056) <= std_logic_vector(output_X8_Y4_gray);
data_out(1071 downto 1064) <= std_logic_vector(output_X8_Y5_gray);
data_out(1079 downto 1072) <= std_logic_vector(output_X8_Y6_gray);
data_out(1087 downto 1080) <= std_logic_vector(output_X8_Y7_gray);
data_out(1095 downto 1088) <= std_logic_vector(output_X8_Y8_gray);
data_out(1103 downto 1096) <= std_logic_vector(output_X8_Y9_gray);
data_out(1111 downto 1104) <= std_logic_vector(output_X8_Y10_gray);
data_out(1119 downto 1112) <= std_logic_vector(output_X8_Y11_gray);
data_out(1127 downto 1120) <= std_logic_vector(output_X8_Y12_gray);
data_out(1135 downto 1128) <= std_logic_vector(output_X8_Y13_gray);
data_out(1143 downto 1136) <= std_logic_vector(output_X8_Y14_gray);
data_out(1151 downto 1144) <= std_logic_vector(output_X8_Y15_gray);
data_out(1159 downto 1152) <= std_logic_vector(output_X9_Y0_gray);
data_out(1167 downto 1160) <= std_logic_vector(output_X9_Y1_gray);
data_out(1175 downto 1168) <= std_logic_vector(output_X9_Y2_gray);
data_out(1183 downto 1176) <= std_logic_vector(output_X9_Y3_gray);
data_out(1191 downto 1184) <= std_logic_vector(output_X9_Y4_gray);
data_out(1199 downto 1192) <= std_logic_vector(output_X9_Y5_gray);
data_out(1207 downto 1200) <= std_logic_vector(output_X9_Y6_gray);
data_out(1215 downto 1208) <= std_logic_vector(output_X9_Y7_gray);
data_out(1223 downto 1216) <= std_logic_vector(output_X9_Y8_gray);
data_out(1231 downto 1224) <= std_logic_vector(output_X9_Y9_gray);
data_out(1239 downto 1232) <= std_logic_vector(output_X9_Y10_gray);
data_out(1247 downto 1240) <= std_logic_vector(output_X9_Y11_gray);
data_out(1255 downto 1248) <= std_logic_vector(output_X9_Y12_gray);
data_out(1263 downto 1256) <= std_logic_vector(output_X9_Y13_gray);
data_out(1271 downto 1264) <= std_logic_vector(output_X9_Y14_gray);
data_out(1279 downto 1272) <= std_logic_vector(output_X9_Y15_gray);
data_out(1287 downto 1280) <= std_logic_vector(output_X10_Y0_gray);
data_out(1295 downto 1288) <= std_logic_vector(output_X10_Y1_gray);
data_out(1303 downto 1296) <= std_logic_vector(output_X10_Y2_gray);
data_out(1311 downto 1304) <= std_logic_vector(output_X10_Y3_gray);
data_out(1319 downto 1312) <= std_logic_vector(output_X10_Y4_gray);
data_out(1327 downto 1320) <= std_logic_vector(output_X10_Y5_gray);
data_out(1335 downto 1328) <= std_logic_vector(output_X10_Y6_gray);
data_out(1343 downto 1336) <= std_logic_vector(output_X10_Y7_gray);
data_out(1351 downto 1344) <= std_logic_vector(output_X10_Y8_gray);
data_out(1359 downto 1352) <= std_logic_vector(output_X10_Y9_gray);
data_out(1367 downto 1360) <= std_logic_vector(output_X10_Y10_gray);
data_out(1375 downto 1368) <= std_logic_vector(output_X10_Y11_gray);
data_out(1383 downto 1376) <= std_logic_vector(output_X10_Y12_gray);
data_out(1391 downto 1384) <= std_logic_vector(output_X10_Y13_gray);
data_out(1399 downto 1392) <= std_logic_vector(output_X10_Y14_gray);
data_out(1407 downto 1400) <= std_logic_vector(output_X10_Y15_gray);
data_out(1415 downto 1408) <= std_logic_vector(output_X11_Y0_gray);
data_out(1423 downto 1416) <= std_logic_vector(output_X11_Y1_gray);
data_out(1431 downto 1424) <= std_logic_vector(output_X11_Y2_gray);
data_out(1439 downto 1432) <= std_logic_vector(output_X11_Y3_gray);
data_out(1447 downto 1440) <= std_logic_vector(output_X11_Y4_gray);
data_out(1455 downto 1448) <= std_logic_vector(output_X11_Y5_gray);
data_out(1463 downto 1456) <= std_logic_vector(output_X11_Y6_gray);
data_out(1471 downto 1464) <= std_logic_vector(output_X11_Y7_gray);
data_out(1479 downto 1472) <= std_logic_vector(output_X11_Y8_gray);
data_out(1487 downto 1480) <= std_logic_vector(output_X11_Y9_gray);
data_out(1495 downto 1488) <= std_logic_vector(output_X11_Y10_gray);
data_out(1503 downto 1496) <= std_logic_vector(output_X11_Y11_gray);
data_out(1511 downto 1504) <= std_logic_vector(output_X11_Y12_gray);
data_out(1519 downto 1512) <= std_logic_vector(output_X11_Y13_gray);
data_out(1527 downto 1520) <= std_logic_vector(output_X11_Y14_gray);
data_out(1535 downto 1528) <= std_logic_vector(output_X11_Y15_gray);
data_out(1543 downto 1536) <= std_logic_vector(output_X12_Y0_gray);
data_out(1551 downto 1544) <= std_logic_vector(output_X12_Y1_gray);
data_out(1559 downto 1552) <= std_logic_vector(output_X12_Y2_gray);
data_out(1567 downto 1560) <= std_logic_vector(output_X12_Y3_gray);
data_out(1575 downto 1568) <= std_logic_vector(output_X12_Y4_gray);
data_out(1583 downto 1576) <= std_logic_vector(output_X12_Y5_gray);
data_out(1591 downto 1584) <= std_logic_vector(output_X12_Y6_gray);
data_out(1599 downto 1592) <= std_logic_vector(output_X12_Y7_gray);
data_out(1607 downto 1600) <= std_logic_vector(output_X12_Y8_gray);
data_out(1615 downto 1608) <= std_logic_vector(output_X12_Y9_gray);
data_out(1623 downto 1616) <= std_logic_vector(output_X12_Y10_gray);
data_out(1631 downto 1624) <= std_logic_vector(output_X12_Y11_gray);
data_out(1639 downto 1632) <= std_logic_vector(output_X12_Y12_gray);
data_out(1647 downto 1640) <= std_logic_vector(output_X12_Y13_gray);
data_out(1655 downto 1648) <= std_logic_vector(output_X12_Y14_gray);
data_out(1663 downto 1656) <= std_logic_vector(output_X12_Y15_gray);
data_out(1671 downto 1664) <= std_logic_vector(output_X13_Y0_gray);
data_out(1679 downto 1672) <= std_logic_vector(output_X13_Y1_gray);
data_out(1687 downto 1680) <= std_logic_vector(output_X13_Y2_gray);
data_out(1695 downto 1688) <= std_logic_vector(output_X13_Y3_gray);
data_out(1703 downto 1696) <= std_logic_vector(output_X13_Y4_gray);
data_out(1711 downto 1704) <= std_logic_vector(output_X13_Y5_gray);
data_out(1719 downto 1712) <= std_logic_vector(output_X13_Y6_gray);
data_out(1727 downto 1720) <= std_logic_vector(output_X13_Y7_gray);
data_out(1735 downto 1728) <= std_logic_vector(output_X13_Y8_gray);
data_out(1743 downto 1736) <= std_logic_vector(output_X13_Y9_gray);
data_out(1751 downto 1744) <= std_logic_vector(output_X13_Y10_gray);
data_out(1759 downto 1752) <= std_logic_vector(output_X13_Y11_gray);
data_out(1767 downto 1760) <= std_logic_vector(output_X13_Y12_gray);
data_out(1775 downto 1768) <= std_logic_vector(output_X13_Y13_gray);
data_out(1783 downto 1776) <= std_logic_vector(output_X13_Y14_gray);
data_out(1791 downto 1784) <= std_logic_vector(output_X13_Y15_gray);
data_out(1799 downto 1792) <= std_logic_vector(output_X14_Y0_gray);
data_out(1807 downto 1800) <= std_logic_vector(output_X14_Y1_gray);
data_out(1815 downto 1808) <= std_logic_vector(output_X14_Y2_gray);
data_out(1823 downto 1816) <= std_logic_vector(output_X14_Y3_gray);
data_out(1831 downto 1824) <= std_logic_vector(output_X14_Y4_gray);
data_out(1839 downto 1832) <= std_logic_vector(output_X14_Y5_gray);
data_out(1847 downto 1840) <= std_logic_vector(output_X14_Y6_gray);
data_out(1855 downto 1848) <= std_logic_vector(output_X14_Y7_gray);
data_out(1863 downto 1856) <= std_logic_vector(output_X14_Y8_gray);
data_out(1871 downto 1864) <= std_logic_vector(output_X14_Y9_gray);
data_out(1879 downto 1872) <= std_logic_vector(output_X14_Y10_gray);
data_out(1887 downto 1880) <= std_logic_vector(output_X14_Y11_gray);
data_out(1895 downto 1888) <= std_logic_vector(output_X14_Y12_gray);
data_out(1903 downto 1896) <= std_logic_vector(output_X14_Y13_gray);
data_out(1911 downto 1904) <= std_logic_vector(output_X14_Y14_gray);
data_out(1919 downto 1912) <= std_logic_vector(output_X14_Y15_gray);
data_out(1927 downto 1920) <= std_logic_vector(output_X15_Y0_gray);
data_out(1935 downto 1928) <= std_logic_vector(output_X15_Y1_gray);
data_out(1943 downto 1936) <= std_logic_vector(output_X15_Y2_gray);
data_out(1951 downto 1944) <= std_logic_vector(output_X15_Y3_gray);
data_out(1959 downto 1952) <= std_logic_vector(output_X15_Y4_gray);
data_out(1967 downto 1960) <= std_logic_vector(output_X15_Y5_gray);
data_out(1975 downto 1968) <= std_logic_vector(output_X15_Y6_gray);
data_out(1983 downto 1976) <= std_logic_vector(output_X15_Y7_gray);
data_out(1991 downto 1984) <= std_logic_vector(output_X15_Y8_gray);
data_out(1999 downto 1992) <= std_logic_vector(output_X15_Y9_gray);
data_out(2007 downto 2000) <= std_logic_vector(output_X15_Y10_gray);
data_out(2015 downto 2008) <= std_logic_vector(output_X15_Y11_gray);
data_out(2023 downto 2016) <= std_logic_vector(output_X15_Y12_gray);
data_out(2031 downto 2024) <= std_logic_vector(output_X15_Y13_gray);
data_out(2039 downto 2032) <= std_logic_vector(output_X15_Y14_gray);
data_out(2047 downto 2040) <= std_logic_vector(output_X15_Y15_gray);



    --      INSERT HERE YOUR VHDL CODE
output_X0_Y0_gray <= input_X0_Y0_r when input_X0_Y0_r >= input_X0_Y0_b and input_X0_Y0_r >= input_X0_Y0_g else input_X0_Y0_g when input_X0_Y0_g >= input_X0_Y0_b else input_X0_Y0_b;
output_X0_Y1_gray <= input_X0_Y1_r when input_X0_Y1_r >= input_X0_Y1_b and input_X0_Y1_r >= input_X0_Y1_g else input_X0_Y1_g when input_X0_Y1_g >= input_X0_Y1_b else input_X0_Y1_b;
output_X0_Y2_gray <= input_X0_Y2_r when input_X0_Y2_r >= input_X0_Y2_b and input_X0_Y2_r >= input_X0_Y2_g else input_X0_Y2_g when input_X0_Y2_g >= input_X0_Y2_b else input_X0_Y2_b;
output_X0_Y3_gray <= input_X0_Y3_r when input_X0_Y3_r >= input_X0_Y3_b and input_X0_Y3_r >= input_X0_Y3_g else input_X0_Y3_g when input_X0_Y3_g >= input_X0_Y3_b else input_X0_Y3_b;
output_X0_Y4_gray <= input_X0_Y4_r when input_X0_Y4_r >= input_X0_Y4_b and input_X0_Y4_r >= input_X0_Y4_g else input_X0_Y4_g when input_X0_Y4_g >= input_X0_Y4_b else input_X0_Y4_b;
output_X0_Y5_gray <= input_X0_Y5_r when input_X0_Y5_r >= input_X0_Y5_b and input_X0_Y5_r >= input_X0_Y5_g else input_X0_Y5_g when input_X0_Y5_g >= input_X0_Y5_b else input_X0_Y5_b;
output_X0_Y6_gray <= input_X0_Y6_r when input_X0_Y6_r >= input_X0_Y6_b and input_X0_Y6_r >= input_X0_Y6_g else input_X0_Y6_g when input_X0_Y6_g >= input_X0_Y6_b else input_X0_Y6_b;
output_X0_Y7_gray <= input_X0_Y7_r when input_X0_Y7_r >= input_X0_Y7_b and input_X0_Y7_r >= input_X0_Y7_g else input_X0_Y7_g when input_X0_Y7_g >= input_X0_Y7_b else input_X0_Y7_b;
output_X0_Y8_gray <= input_X0_Y8_r when input_X0_Y8_r >= input_X0_Y8_b and input_X0_Y8_r >= input_X0_Y8_g else input_X0_Y8_g when input_X0_Y8_g >= input_X0_Y8_b else input_X0_Y8_b;
output_X0_Y9_gray <= input_X0_Y9_r when input_X0_Y9_r >= input_X0_Y9_b and input_X0_Y9_r >= input_X0_Y9_g else input_X0_Y9_g when input_X0_Y9_g >= input_X0_Y9_b else input_X0_Y9_b;
output_X0_Y10_gray <= input_X0_Y10_r when input_X0_Y10_r >= input_X0_Y10_b and input_X0_Y10_r >= input_X0_Y10_g else input_X0_Y10_g when input_X0_Y10_g >= input_X0_Y10_b else input_X0_Y10_b;
output_X0_Y11_gray <= input_X0_Y11_r when input_X0_Y11_r >= input_X0_Y11_b and input_X0_Y11_r >= input_X0_Y11_g else input_X0_Y11_g when input_X0_Y11_g >= input_X0_Y11_b else input_X0_Y11_b;
output_X0_Y12_gray <= input_X0_Y12_r when input_X0_Y12_r >= input_X0_Y12_b and input_X0_Y12_r >= input_X0_Y12_g else input_X0_Y12_g when input_X0_Y12_g >= input_X0_Y12_b else input_X0_Y12_b;
output_X0_Y13_gray <= input_X0_Y13_r when input_X0_Y13_r >= input_X0_Y13_b and input_X0_Y13_r >= input_X0_Y13_g else input_X0_Y13_g when input_X0_Y13_g >= input_X0_Y13_b else input_X0_Y13_b;
output_X0_Y14_gray <= input_X0_Y14_r when input_X0_Y14_r >= input_X0_Y14_b and input_X0_Y14_r >= input_X0_Y14_g else input_X0_Y14_g when input_X0_Y14_g >= input_X0_Y14_b else input_X0_Y14_b;
output_X0_Y15_gray <= input_X0_Y15_r when input_X0_Y15_r >= input_X0_Y15_b and input_X0_Y15_r >= input_X0_Y15_g else input_X0_Y15_g when input_X0_Y15_g >= input_X0_Y15_b else input_X0_Y15_b;
output_X1_Y0_gray <= input_X1_Y0_r when input_X1_Y0_r >= input_X1_Y0_b and input_X1_Y0_r >= input_X1_Y0_g else input_X1_Y0_g when input_X1_Y0_g >= input_X1_Y0_b else input_X1_Y0_b;
output_X1_Y1_gray <= input_X1_Y1_r when input_X1_Y1_r >= input_X1_Y1_b and input_X1_Y1_r >= input_X1_Y1_g else input_X1_Y1_g when input_X1_Y1_g >= input_X1_Y1_b else input_X1_Y1_b;
output_X1_Y2_gray <= input_X1_Y2_r when input_X1_Y2_r >= input_X1_Y2_b and input_X1_Y2_r >= input_X1_Y2_g else input_X1_Y2_g when input_X1_Y2_g >= input_X1_Y2_b else input_X1_Y2_b;
output_X1_Y3_gray <= input_X1_Y3_r when input_X1_Y3_r >= input_X1_Y3_b and input_X1_Y3_r >= input_X1_Y3_g else input_X1_Y3_g when input_X1_Y3_g >= input_X1_Y3_b else input_X1_Y3_b;
output_X1_Y4_gray <= input_X1_Y4_r when input_X1_Y4_r >= input_X1_Y4_b and input_X1_Y4_r >= input_X1_Y4_g else input_X1_Y4_g when input_X1_Y4_g >= input_X1_Y4_b else input_X1_Y4_b;
output_X1_Y5_gray <= input_X1_Y5_r when input_X1_Y5_r >= input_X1_Y5_b and input_X1_Y5_r >= input_X1_Y5_g else input_X1_Y5_g when input_X1_Y5_g >= input_X1_Y5_b else input_X1_Y5_b;
output_X1_Y6_gray <= input_X1_Y6_r when input_X1_Y6_r >= input_X1_Y6_b and input_X1_Y6_r >= input_X1_Y6_g else input_X1_Y6_g when input_X1_Y6_g >= input_X1_Y6_b else input_X1_Y6_b;
output_X1_Y7_gray <= input_X1_Y7_r when input_X1_Y7_r >= input_X1_Y7_b and input_X1_Y7_r >= input_X1_Y7_g else input_X1_Y7_g when input_X1_Y7_g >= input_X1_Y7_b else input_X1_Y7_b;
output_X1_Y8_gray <= input_X1_Y8_r when input_X1_Y8_r >= input_X1_Y8_b and input_X1_Y8_r >= input_X1_Y8_g else input_X1_Y8_g when input_X1_Y8_g >= input_X1_Y8_b else input_X1_Y8_b;
output_X1_Y9_gray <= input_X1_Y9_r when input_X1_Y9_r >= input_X1_Y9_b and input_X1_Y9_r >= input_X1_Y9_g else input_X1_Y9_g when input_X1_Y9_g >= input_X1_Y9_b else input_X1_Y9_b;
output_X1_Y10_gray <= input_X1_Y10_r when input_X1_Y10_r >= input_X1_Y10_b and input_X1_Y10_r >= input_X1_Y10_g else input_X1_Y10_g when input_X1_Y10_g >= input_X1_Y10_b else input_X1_Y10_b;
output_X1_Y11_gray <= input_X1_Y11_r when input_X1_Y11_r >= input_X1_Y11_b and input_X1_Y11_r >= input_X1_Y11_g else input_X1_Y11_g when input_X1_Y11_g >= input_X1_Y11_b else input_X1_Y11_b;
output_X1_Y12_gray <= input_X1_Y12_r when input_X1_Y12_r >= input_X1_Y12_b and input_X1_Y12_r >= input_X1_Y12_g else input_X1_Y12_g when input_X1_Y12_g >= input_X1_Y12_b else input_X1_Y12_b;
output_X1_Y13_gray <= input_X1_Y13_r when input_X1_Y13_r >= input_X1_Y13_b and input_X1_Y13_r >= input_X1_Y13_g else input_X1_Y13_g when input_X1_Y13_g >= input_X1_Y13_b else input_X1_Y13_b;
output_X1_Y14_gray <= input_X1_Y14_r when input_X1_Y14_r >= input_X1_Y14_b and input_X1_Y14_r >= input_X1_Y14_g else input_X1_Y14_g when input_X1_Y14_g >= input_X1_Y14_b else input_X1_Y14_b;
output_X1_Y15_gray <= input_X1_Y15_r when input_X1_Y15_r >= input_X1_Y15_b and input_X1_Y15_r >= input_X1_Y15_g else input_X1_Y15_g when input_X1_Y15_g >= input_X1_Y15_b else input_X1_Y15_b;
output_X2_Y0_gray <= input_X2_Y0_r when input_X2_Y0_r >= input_X2_Y0_b and input_X2_Y0_r >= input_X2_Y0_g else input_X2_Y0_g when input_X2_Y0_g >= input_X2_Y0_b else input_X2_Y0_b;
output_X2_Y1_gray <= input_X2_Y1_r when input_X2_Y1_r >= input_X2_Y1_b and input_X2_Y1_r >= input_X2_Y1_g else input_X2_Y1_g when input_X2_Y1_g >= input_X2_Y1_b else input_X2_Y1_b;
output_X2_Y2_gray <= input_X2_Y2_r when input_X2_Y2_r >= input_X2_Y2_b and input_X2_Y2_r >= input_X2_Y2_g else input_X2_Y2_g when input_X2_Y2_g >= input_X2_Y2_b else input_X2_Y2_b;
output_X2_Y3_gray <= input_X2_Y3_r when input_X2_Y3_r >= input_X2_Y3_b and input_X2_Y3_r >= input_X2_Y3_g else input_X2_Y3_g when input_X2_Y3_g >= input_X2_Y3_b else input_X2_Y3_b;
output_X2_Y4_gray <= input_X2_Y4_r when input_X2_Y4_r >= input_X2_Y4_b and input_X2_Y4_r >= input_X2_Y4_g else input_X2_Y4_g when input_X2_Y4_g >= input_X2_Y4_b else input_X2_Y4_b;
output_X2_Y5_gray <= input_X2_Y5_r when input_X2_Y5_r >= input_X2_Y5_b and input_X2_Y5_r >= input_X2_Y5_g else input_X2_Y5_g when input_X2_Y5_g >= input_X2_Y5_b else input_X2_Y5_b;
output_X2_Y6_gray <= input_X2_Y6_r when input_X2_Y6_r >= input_X2_Y6_b and input_X2_Y6_r >= input_X2_Y6_g else input_X2_Y6_g when input_X2_Y6_g >= input_X2_Y6_b else input_X2_Y6_b;
output_X2_Y7_gray <= input_X2_Y7_r when input_X2_Y7_r >= input_X2_Y7_b and input_X2_Y7_r >= input_X2_Y7_g else input_X2_Y7_g when input_X2_Y7_g >= input_X2_Y7_b else input_X2_Y7_b;
output_X2_Y8_gray <= input_X2_Y8_r when input_X2_Y8_r >= input_X2_Y8_b and input_X2_Y8_r >= input_X2_Y8_g else input_X2_Y8_g when input_X2_Y8_g >= input_X2_Y8_b else input_X2_Y8_b;
output_X2_Y9_gray <= input_X2_Y9_r when input_X2_Y9_r >= input_X2_Y9_b and input_X2_Y9_r >= input_X2_Y9_g else input_X2_Y9_g when input_X2_Y9_g >= input_X2_Y9_b else input_X2_Y9_b;
output_X2_Y10_gray <= input_X2_Y10_r when input_X2_Y10_r >= input_X2_Y10_b and input_X2_Y10_r >= input_X2_Y10_g else input_X2_Y10_g when input_X2_Y10_g >= input_X2_Y10_b else input_X2_Y10_b;
output_X2_Y11_gray <= input_X2_Y11_r when input_X2_Y11_r >= input_X2_Y11_b and input_X2_Y11_r >= input_X2_Y11_g else input_X2_Y11_g when input_X2_Y11_g >= input_X2_Y11_b else input_X2_Y11_b;
output_X2_Y12_gray <= input_X2_Y12_r when input_X2_Y12_r >= input_X2_Y12_b and input_X2_Y12_r >= input_X2_Y12_g else input_X2_Y12_g when input_X2_Y12_g >= input_X2_Y12_b else input_X2_Y12_b;
output_X2_Y13_gray <= input_X2_Y13_r when input_X2_Y13_r >= input_X2_Y13_b and input_X2_Y13_r >= input_X2_Y13_g else input_X2_Y13_g when input_X2_Y13_g >= input_X2_Y13_b else input_X2_Y13_b;
output_X2_Y14_gray <= input_X2_Y14_r when input_X2_Y14_r >= input_X2_Y14_b and input_X2_Y14_r >= input_X2_Y14_g else input_X2_Y14_g when input_X2_Y14_g >= input_X2_Y14_b else input_X2_Y14_b;
output_X2_Y15_gray <= input_X2_Y15_r when input_X2_Y15_r >= input_X2_Y15_b and input_X2_Y15_r >= input_X2_Y15_g else input_X2_Y15_g when input_X2_Y15_g >= input_X2_Y15_b else input_X2_Y15_b;
output_X3_Y0_gray <= input_X3_Y0_r when input_X3_Y0_r >= input_X3_Y0_b and input_X3_Y0_r >= input_X3_Y0_g else input_X3_Y0_g when input_X3_Y0_g >= input_X3_Y0_b else input_X3_Y0_b;
output_X3_Y1_gray <= input_X3_Y1_r when input_X3_Y1_r >= input_X3_Y1_b and input_X3_Y1_r >= input_X3_Y1_g else input_X3_Y1_g when input_X3_Y1_g >= input_X3_Y1_b else input_X3_Y1_b;
output_X3_Y2_gray <= input_X3_Y2_r when input_X3_Y2_r >= input_X3_Y2_b and input_X3_Y2_r >= input_X3_Y2_g else input_X3_Y2_g when input_X3_Y2_g >= input_X3_Y2_b else input_X3_Y2_b;
output_X3_Y3_gray <= input_X3_Y3_r when input_X3_Y3_r >= input_X3_Y3_b and input_X3_Y3_r >= input_X3_Y3_g else input_X3_Y3_g when input_X3_Y3_g >= input_X3_Y3_b else input_X3_Y3_b;
output_X3_Y4_gray <= input_X3_Y4_r when input_X3_Y4_r >= input_X3_Y4_b and input_X3_Y4_r >= input_X3_Y4_g else input_X3_Y4_g when input_X3_Y4_g >= input_X3_Y4_b else input_X3_Y4_b;
output_X3_Y5_gray <= input_X3_Y5_r when input_X3_Y5_r >= input_X3_Y5_b and input_X3_Y5_r >= input_X3_Y5_g else input_X3_Y5_g when input_X3_Y5_g >= input_X3_Y5_b else input_X3_Y5_b;
output_X3_Y6_gray <= input_X3_Y6_r when input_X3_Y6_r >= input_X3_Y6_b and input_X3_Y6_r >= input_X3_Y6_g else input_X3_Y6_g when input_X3_Y6_g >= input_X3_Y6_b else input_X3_Y6_b;
output_X3_Y7_gray <= input_X3_Y7_r when input_X3_Y7_r >= input_X3_Y7_b and input_X3_Y7_r >= input_X3_Y7_g else input_X3_Y7_g when input_X3_Y7_g >= input_X3_Y7_b else input_X3_Y7_b;
output_X3_Y8_gray <= input_X3_Y8_r when input_X3_Y8_r >= input_X3_Y8_b and input_X3_Y8_r >= input_X3_Y8_g else input_X3_Y8_g when input_X3_Y8_g >= input_X3_Y8_b else input_X3_Y8_b;
output_X3_Y9_gray <= input_X3_Y9_r when input_X3_Y9_r >= input_X3_Y9_b and input_X3_Y9_r >= input_X3_Y9_g else input_X3_Y9_g when input_X3_Y9_g >= input_X3_Y9_b else input_X3_Y9_b;
output_X3_Y10_gray <= input_X3_Y10_r when input_X3_Y10_r >= input_X3_Y10_b and input_X3_Y10_r >= input_X3_Y10_g else input_X3_Y10_g when input_X3_Y10_g >= input_X3_Y10_b else input_X3_Y10_b;
output_X3_Y11_gray <= input_X3_Y11_r when input_X3_Y11_r >= input_X3_Y11_b and input_X3_Y11_r >= input_X3_Y11_g else input_X3_Y11_g when input_X3_Y11_g >= input_X3_Y11_b else input_X3_Y11_b;
output_X3_Y12_gray <= input_X3_Y12_r when input_X3_Y12_r >= input_X3_Y12_b and input_X3_Y12_r >= input_X3_Y12_g else input_X3_Y12_g when input_X3_Y12_g >= input_X3_Y12_b else input_X3_Y12_b;
output_X3_Y13_gray <= input_X3_Y13_r when input_X3_Y13_r >= input_X3_Y13_b and input_X3_Y13_r >= input_X3_Y13_g else input_X3_Y13_g when input_X3_Y13_g >= input_X3_Y13_b else input_X3_Y13_b;
output_X3_Y14_gray <= input_X3_Y14_r when input_X3_Y14_r >= input_X3_Y14_b and input_X3_Y14_r >= input_X3_Y14_g else input_X3_Y14_g when input_X3_Y14_g >= input_X3_Y14_b else input_X3_Y14_b;
output_X3_Y15_gray <= input_X3_Y15_r when input_X3_Y15_r >= input_X3_Y15_b and input_X3_Y15_r >= input_X3_Y15_g else input_X3_Y15_g when input_X3_Y15_g >= input_X3_Y15_b else input_X3_Y15_b;
output_X4_Y0_gray <= input_X4_Y0_r when input_X4_Y0_r >= input_X4_Y0_b and input_X4_Y0_r >= input_X4_Y0_g else input_X4_Y0_g when input_X4_Y0_g >= input_X4_Y0_b else input_X4_Y0_b;
output_X4_Y1_gray <= input_X4_Y1_r when input_X4_Y1_r >= input_X4_Y1_b and input_X4_Y1_r >= input_X4_Y1_g else input_X4_Y1_g when input_X4_Y1_g >= input_X4_Y1_b else input_X4_Y1_b;
output_X4_Y2_gray <= input_X4_Y2_r when input_X4_Y2_r >= input_X4_Y2_b and input_X4_Y2_r >= input_X4_Y2_g else input_X4_Y2_g when input_X4_Y2_g >= input_X4_Y2_b else input_X4_Y2_b;
output_X4_Y3_gray <= input_X4_Y3_r when input_X4_Y3_r >= input_X4_Y3_b and input_X4_Y3_r >= input_X4_Y3_g else input_X4_Y3_g when input_X4_Y3_g >= input_X4_Y3_b else input_X4_Y3_b;
output_X4_Y4_gray <= input_X4_Y4_r when input_X4_Y4_r >= input_X4_Y4_b and input_X4_Y4_r >= input_X4_Y4_g else input_X4_Y4_g when input_X4_Y4_g >= input_X4_Y4_b else input_X4_Y4_b;
output_X4_Y5_gray <= input_X4_Y5_r when input_X4_Y5_r >= input_X4_Y5_b and input_X4_Y5_r >= input_X4_Y5_g else input_X4_Y5_g when input_X4_Y5_g >= input_X4_Y5_b else input_X4_Y5_b;
output_X4_Y6_gray <= input_X4_Y6_r when input_X4_Y6_r >= input_X4_Y6_b and input_X4_Y6_r >= input_X4_Y6_g else input_X4_Y6_g when input_X4_Y6_g >= input_X4_Y6_b else input_X4_Y6_b;
output_X4_Y7_gray <= input_X4_Y7_r when input_X4_Y7_r >= input_X4_Y7_b and input_X4_Y7_r >= input_X4_Y7_g else input_X4_Y7_g when input_X4_Y7_g >= input_X4_Y7_b else input_X4_Y7_b;
output_X4_Y8_gray <= input_X4_Y8_r when input_X4_Y8_r >= input_X4_Y8_b and input_X4_Y8_r >= input_X4_Y8_g else input_X4_Y8_g when input_X4_Y8_g >= input_X4_Y8_b else input_X4_Y8_b;
output_X4_Y9_gray <= input_X4_Y9_r when input_X4_Y9_r >= input_X4_Y9_b and input_X4_Y9_r >= input_X4_Y9_g else input_X4_Y9_g when input_X4_Y9_g >= input_X4_Y9_b else input_X4_Y9_b;
output_X4_Y10_gray <= input_X4_Y10_r when input_X4_Y10_r >= input_X4_Y10_b and input_X4_Y10_r >= input_X4_Y10_g else input_X4_Y10_g when input_X4_Y10_g >= input_X4_Y10_b else input_X4_Y10_b;
output_X4_Y11_gray <= input_X4_Y11_r when input_X4_Y11_r >= input_X4_Y11_b and input_X4_Y11_r >= input_X4_Y11_g else input_X4_Y11_g when input_X4_Y11_g >= input_X4_Y11_b else input_X4_Y11_b;
output_X4_Y12_gray <= input_X4_Y12_r when input_X4_Y12_r >= input_X4_Y12_b and input_X4_Y12_r >= input_X4_Y12_g else input_X4_Y12_g when input_X4_Y12_g >= input_X4_Y12_b else input_X4_Y12_b;
output_X4_Y13_gray <= input_X4_Y13_r when input_X4_Y13_r >= input_X4_Y13_b and input_X4_Y13_r >= input_X4_Y13_g else input_X4_Y13_g when input_X4_Y13_g >= input_X4_Y13_b else input_X4_Y13_b;
output_X4_Y14_gray <= input_X4_Y14_r when input_X4_Y14_r >= input_X4_Y14_b and input_X4_Y14_r >= input_X4_Y14_g else input_X4_Y14_g when input_X4_Y14_g >= input_X4_Y14_b else input_X4_Y14_b;
output_X4_Y15_gray <= input_X4_Y15_r when input_X4_Y15_r >= input_X4_Y15_b and input_X4_Y15_r >= input_X4_Y15_g else input_X4_Y15_g when input_X4_Y15_g >= input_X4_Y15_b else input_X4_Y15_b;
output_X5_Y0_gray <= input_X5_Y0_r when input_X5_Y0_r >= input_X5_Y0_b and input_X5_Y0_r >= input_X5_Y0_g else input_X5_Y0_g when input_X5_Y0_g >= input_X5_Y0_b else input_X5_Y0_b;
output_X5_Y1_gray <= input_X5_Y1_r when input_X5_Y1_r >= input_X5_Y1_b and input_X5_Y1_r >= input_X5_Y1_g else input_X5_Y1_g when input_X5_Y1_g >= input_X5_Y1_b else input_X5_Y1_b;
output_X5_Y2_gray <= input_X5_Y2_r when input_X5_Y2_r >= input_X5_Y2_b and input_X5_Y2_r >= input_X5_Y2_g else input_X5_Y2_g when input_X5_Y2_g >= input_X5_Y2_b else input_X5_Y2_b;
output_X5_Y3_gray <= input_X5_Y3_r when input_X5_Y3_r >= input_X5_Y3_b and input_X5_Y3_r >= input_X5_Y3_g else input_X5_Y3_g when input_X5_Y3_g >= input_X5_Y3_b else input_X5_Y3_b;
output_X5_Y4_gray <= input_X5_Y4_r when input_X5_Y4_r >= input_X5_Y4_b and input_X5_Y4_r >= input_X5_Y4_g else input_X5_Y4_g when input_X5_Y4_g >= input_X5_Y4_b else input_X5_Y4_b;
output_X5_Y5_gray <= input_X5_Y5_r when input_X5_Y5_r >= input_X5_Y5_b and input_X5_Y5_r >= input_X5_Y5_g else input_X5_Y5_g when input_X5_Y5_g >= input_X5_Y5_b else input_X5_Y5_b;
output_X5_Y6_gray <= input_X5_Y6_r when input_X5_Y6_r >= input_X5_Y6_b and input_X5_Y6_r >= input_X5_Y6_g else input_X5_Y6_g when input_X5_Y6_g >= input_X5_Y6_b else input_X5_Y6_b;
output_X5_Y7_gray <= input_X5_Y7_r when input_X5_Y7_r >= input_X5_Y7_b and input_X5_Y7_r >= input_X5_Y7_g else input_X5_Y7_g when input_X5_Y7_g >= input_X5_Y7_b else input_X5_Y7_b;
output_X5_Y8_gray <= input_X5_Y8_r when input_X5_Y8_r >= input_X5_Y8_b and input_X5_Y8_r >= input_X5_Y8_g else input_X5_Y8_g when input_X5_Y8_g >= input_X5_Y8_b else input_X5_Y8_b;
output_X5_Y9_gray <= input_X5_Y9_r when input_X5_Y9_r >= input_X5_Y9_b and input_X5_Y9_r >= input_X5_Y9_g else input_X5_Y9_g when input_X5_Y9_g >= input_X5_Y9_b else input_X5_Y9_b;
output_X5_Y10_gray <= input_X5_Y10_r when input_X5_Y10_r >= input_X5_Y10_b and input_X5_Y10_r >= input_X5_Y10_g else input_X5_Y10_g when input_X5_Y10_g >= input_X5_Y10_b else input_X5_Y10_b;
output_X5_Y11_gray <= input_X5_Y11_r when input_X5_Y11_r >= input_X5_Y11_b and input_X5_Y11_r >= input_X5_Y11_g else input_X5_Y11_g when input_X5_Y11_g >= input_X5_Y11_b else input_X5_Y11_b;
output_X5_Y12_gray <= input_X5_Y12_r when input_X5_Y12_r >= input_X5_Y12_b and input_X5_Y12_r >= input_X5_Y12_g else input_X5_Y12_g when input_X5_Y12_g >= input_X5_Y12_b else input_X5_Y12_b;
output_X5_Y13_gray <= input_X5_Y13_r when input_X5_Y13_r >= input_X5_Y13_b and input_X5_Y13_r >= input_X5_Y13_g else input_X5_Y13_g when input_X5_Y13_g >= input_X5_Y13_b else input_X5_Y13_b;
output_X5_Y14_gray <= input_X5_Y14_r when input_X5_Y14_r >= input_X5_Y14_b and input_X5_Y14_r >= input_X5_Y14_g else input_X5_Y14_g when input_X5_Y14_g >= input_X5_Y14_b else input_X5_Y14_b;
output_X5_Y15_gray <= input_X5_Y15_r when input_X5_Y15_r >= input_X5_Y15_b and input_X5_Y15_r >= input_X5_Y15_g else input_X5_Y15_g when input_X5_Y15_g >= input_X5_Y15_b else input_X5_Y15_b;
output_X6_Y0_gray <= input_X6_Y0_r when input_X6_Y0_r >= input_X6_Y0_b and input_X6_Y0_r >= input_X6_Y0_g else input_X6_Y0_g when input_X6_Y0_g >= input_X6_Y0_b else input_X6_Y0_b;
output_X6_Y1_gray <= input_X6_Y1_r when input_X6_Y1_r >= input_X6_Y1_b and input_X6_Y1_r >= input_X6_Y1_g else input_X6_Y1_g when input_X6_Y1_g >= input_X6_Y1_b else input_X6_Y1_b;
output_X6_Y2_gray <= input_X6_Y2_r when input_X6_Y2_r >= input_X6_Y2_b and input_X6_Y2_r >= input_X6_Y2_g else input_X6_Y2_g when input_X6_Y2_g >= input_X6_Y2_b else input_X6_Y2_b;
output_X6_Y3_gray <= input_X6_Y3_r when input_X6_Y3_r >= input_X6_Y3_b and input_X6_Y3_r >= input_X6_Y3_g else input_X6_Y3_g when input_X6_Y3_g >= input_X6_Y3_b else input_X6_Y3_b;
output_X6_Y4_gray <= input_X6_Y4_r when input_X6_Y4_r >= input_X6_Y4_b and input_X6_Y4_r >= input_X6_Y4_g else input_X6_Y4_g when input_X6_Y4_g >= input_X6_Y4_b else input_X6_Y4_b;
output_X6_Y5_gray <= input_X6_Y5_r when input_X6_Y5_r >= input_X6_Y5_b and input_X6_Y5_r >= input_X6_Y5_g else input_X6_Y5_g when input_X6_Y5_g >= input_X6_Y5_b else input_X6_Y5_b;
output_X6_Y6_gray <= input_X6_Y6_r when input_X6_Y6_r >= input_X6_Y6_b and input_X6_Y6_r >= input_X6_Y6_g else input_X6_Y6_g when input_X6_Y6_g >= input_X6_Y6_b else input_X6_Y6_b;
output_X6_Y7_gray <= input_X6_Y7_r when input_X6_Y7_r >= input_X6_Y7_b and input_X6_Y7_r >= input_X6_Y7_g else input_X6_Y7_g when input_X6_Y7_g >= input_X6_Y7_b else input_X6_Y7_b;
output_X6_Y8_gray <= input_X6_Y8_r when input_X6_Y8_r >= input_X6_Y8_b and input_X6_Y8_r >= input_X6_Y8_g else input_X6_Y8_g when input_X6_Y8_g >= input_X6_Y8_b else input_X6_Y8_b;
output_X6_Y9_gray <= input_X6_Y9_r when input_X6_Y9_r >= input_X6_Y9_b and input_X6_Y9_r >= input_X6_Y9_g else input_X6_Y9_g when input_X6_Y9_g >= input_X6_Y9_b else input_X6_Y9_b;
output_X6_Y10_gray <= input_X6_Y10_r when input_X6_Y10_r >= input_X6_Y10_b and input_X6_Y10_r >= input_X6_Y10_g else input_X6_Y10_g when input_X6_Y10_g >= input_X6_Y10_b else input_X6_Y10_b;
output_X6_Y11_gray <= input_X6_Y11_r when input_X6_Y11_r >= input_X6_Y11_b and input_X6_Y11_r >= input_X6_Y11_g else input_X6_Y11_g when input_X6_Y11_g >= input_X6_Y11_b else input_X6_Y11_b;
output_X6_Y12_gray <= input_X6_Y12_r when input_X6_Y12_r >= input_X6_Y12_b and input_X6_Y12_r >= input_X6_Y12_g else input_X6_Y12_g when input_X6_Y12_g >= input_X6_Y12_b else input_X6_Y12_b;
output_X6_Y13_gray <= input_X6_Y13_r when input_X6_Y13_r >= input_X6_Y13_b and input_X6_Y13_r >= input_X6_Y13_g else input_X6_Y13_g when input_X6_Y13_g >= input_X6_Y13_b else input_X6_Y13_b;
output_X6_Y14_gray <= input_X6_Y14_r when input_X6_Y14_r >= input_X6_Y14_b and input_X6_Y14_r >= input_X6_Y14_g else input_X6_Y14_g when input_X6_Y14_g >= input_X6_Y14_b else input_X6_Y14_b;
output_X6_Y15_gray <= input_X6_Y15_r when input_X6_Y15_r >= input_X6_Y15_b and input_X6_Y15_r >= input_X6_Y15_g else input_X6_Y15_g when input_X6_Y15_g >= input_X6_Y15_b else input_X6_Y15_b;
output_X7_Y0_gray <= input_X7_Y0_r when input_X7_Y0_r >= input_X7_Y0_b and input_X7_Y0_r >= input_X7_Y0_g else input_X7_Y0_g when input_X7_Y0_g >= input_X7_Y0_b else input_X7_Y0_b;
output_X7_Y1_gray <= input_X7_Y1_r when input_X7_Y1_r >= input_X7_Y1_b and input_X7_Y1_r >= input_X7_Y1_g else input_X7_Y1_g when input_X7_Y1_g >= input_X7_Y1_b else input_X7_Y1_b;
output_X7_Y2_gray <= input_X7_Y2_r when input_X7_Y2_r >= input_X7_Y2_b and input_X7_Y2_r >= input_X7_Y2_g else input_X7_Y2_g when input_X7_Y2_g >= input_X7_Y2_b else input_X7_Y2_b;
output_X7_Y3_gray <= input_X7_Y3_r when input_X7_Y3_r >= input_X7_Y3_b and input_X7_Y3_r >= input_X7_Y3_g else input_X7_Y3_g when input_X7_Y3_g >= input_X7_Y3_b else input_X7_Y3_b;
output_X7_Y4_gray <= input_X7_Y4_r when input_X7_Y4_r >= input_X7_Y4_b and input_X7_Y4_r >= input_X7_Y4_g else input_X7_Y4_g when input_X7_Y4_g >= input_X7_Y4_b else input_X7_Y4_b;
output_X7_Y5_gray <= input_X7_Y5_r when input_X7_Y5_r >= input_X7_Y5_b and input_X7_Y5_r >= input_X7_Y5_g else input_X7_Y5_g when input_X7_Y5_g >= input_X7_Y5_b else input_X7_Y5_b;
output_X7_Y6_gray <= input_X7_Y6_r when input_X7_Y6_r >= input_X7_Y6_b and input_X7_Y6_r >= input_X7_Y6_g else input_X7_Y6_g when input_X7_Y6_g >= input_X7_Y6_b else input_X7_Y6_b;
output_X7_Y7_gray <= input_X7_Y7_r when input_X7_Y7_r >= input_X7_Y7_b and input_X7_Y7_r >= input_X7_Y7_g else input_X7_Y7_g when input_X7_Y7_g >= input_X7_Y7_b else input_X7_Y7_b;
output_X7_Y8_gray <= input_X7_Y8_r when input_X7_Y8_r >= input_X7_Y8_b and input_X7_Y8_r >= input_X7_Y8_g else input_X7_Y8_g when input_X7_Y8_g >= input_X7_Y8_b else input_X7_Y8_b;
output_X7_Y9_gray <= input_X7_Y9_r when input_X7_Y9_r >= input_X7_Y9_b and input_X7_Y9_r >= input_X7_Y9_g else input_X7_Y9_g when input_X7_Y9_g >= input_X7_Y9_b else input_X7_Y9_b;
output_X7_Y10_gray <= input_X7_Y10_r when input_X7_Y10_r >= input_X7_Y10_b and input_X7_Y10_r >= input_X7_Y10_g else input_X7_Y10_g when input_X7_Y10_g >= input_X7_Y10_b else input_X7_Y10_b;
output_X7_Y11_gray <= input_X7_Y11_r when input_X7_Y11_r >= input_X7_Y11_b and input_X7_Y11_r >= input_X7_Y11_g else input_X7_Y11_g when input_X7_Y11_g >= input_X7_Y11_b else input_X7_Y11_b;
output_X7_Y12_gray <= input_X7_Y12_r when input_X7_Y12_r >= input_X7_Y12_b and input_X7_Y12_r >= input_X7_Y12_g else input_X7_Y12_g when input_X7_Y12_g >= input_X7_Y12_b else input_X7_Y12_b;
output_X7_Y13_gray <= input_X7_Y13_r when input_X7_Y13_r >= input_X7_Y13_b and input_X7_Y13_r >= input_X7_Y13_g else input_X7_Y13_g when input_X7_Y13_g >= input_X7_Y13_b else input_X7_Y13_b;
output_X7_Y14_gray <= input_X7_Y14_r when input_X7_Y14_r >= input_X7_Y14_b and input_X7_Y14_r >= input_X7_Y14_g else input_X7_Y14_g when input_X7_Y14_g >= input_X7_Y14_b else input_X7_Y14_b;
output_X7_Y15_gray <= input_X7_Y15_r when input_X7_Y15_r >= input_X7_Y15_b and input_X7_Y15_r >= input_X7_Y15_g else input_X7_Y15_g when input_X7_Y15_g >= input_X7_Y15_b else input_X7_Y15_b;
output_X8_Y0_gray <= input_X8_Y0_r when input_X8_Y0_r >= input_X8_Y0_b and input_X8_Y0_r >= input_X8_Y0_g else input_X8_Y0_g when input_X8_Y0_g >= input_X8_Y0_b else input_X8_Y0_b;
output_X8_Y1_gray <= input_X8_Y1_r when input_X8_Y1_r >= input_X8_Y1_b and input_X8_Y1_r >= input_X8_Y1_g else input_X8_Y1_g when input_X8_Y1_g >= input_X8_Y1_b else input_X8_Y1_b;
output_X8_Y2_gray <= input_X8_Y2_r when input_X8_Y2_r >= input_X8_Y2_b and input_X8_Y2_r >= input_X8_Y2_g else input_X8_Y2_g when input_X8_Y2_g >= input_X8_Y2_b else input_X8_Y2_b;
output_X8_Y3_gray <= input_X8_Y3_r when input_X8_Y3_r >= input_X8_Y3_b and input_X8_Y3_r >= input_X8_Y3_g else input_X8_Y3_g when input_X8_Y3_g >= input_X8_Y3_b else input_X8_Y3_b;
output_X8_Y4_gray <= input_X8_Y4_r when input_X8_Y4_r >= input_X8_Y4_b and input_X8_Y4_r >= input_X8_Y4_g else input_X8_Y4_g when input_X8_Y4_g >= input_X8_Y4_b else input_X8_Y4_b;
output_X8_Y5_gray <= input_X8_Y5_r when input_X8_Y5_r >= input_X8_Y5_b and input_X8_Y5_r >= input_X8_Y5_g else input_X8_Y5_g when input_X8_Y5_g >= input_X8_Y5_b else input_X8_Y5_b;
output_X8_Y6_gray <= input_X8_Y6_r when input_X8_Y6_r >= input_X8_Y6_b and input_X8_Y6_r >= input_X8_Y6_g else input_X8_Y6_g when input_X8_Y6_g >= input_X8_Y6_b else input_X8_Y6_b;
output_X8_Y7_gray <= input_X8_Y7_r when input_X8_Y7_r >= input_X8_Y7_b and input_X8_Y7_r >= input_X8_Y7_g else input_X8_Y7_g when input_X8_Y7_g >= input_X8_Y7_b else input_X8_Y7_b;
output_X8_Y8_gray <= input_X8_Y8_r when input_X8_Y8_r >= input_X8_Y8_b and input_X8_Y8_r >= input_X8_Y8_g else input_X8_Y8_g when input_X8_Y8_g >= input_X8_Y8_b else input_X8_Y8_b;
output_X8_Y9_gray <= input_X8_Y9_r when input_X8_Y9_r >= input_X8_Y9_b and input_X8_Y9_r >= input_X8_Y9_g else input_X8_Y9_g when input_X8_Y9_g >= input_X8_Y9_b else input_X8_Y9_b;
output_X8_Y10_gray <= input_X8_Y10_r when input_X8_Y10_r >= input_X8_Y10_b and input_X8_Y10_r >= input_X8_Y10_g else input_X8_Y10_g when input_X8_Y10_g >= input_X8_Y10_b else input_X8_Y10_b;
output_X8_Y11_gray <= input_X8_Y11_r when input_X8_Y11_r >= input_X8_Y11_b and input_X8_Y11_r >= input_X8_Y11_g else input_X8_Y11_g when input_X8_Y11_g >= input_X8_Y11_b else input_X8_Y11_b;
output_X8_Y12_gray <= input_X8_Y12_r when input_X8_Y12_r >= input_X8_Y12_b and input_X8_Y12_r >= input_X8_Y12_g else input_X8_Y12_g when input_X8_Y12_g >= input_X8_Y12_b else input_X8_Y12_b;
output_X8_Y13_gray <= input_X8_Y13_r when input_X8_Y13_r >= input_X8_Y13_b and input_X8_Y13_r >= input_X8_Y13_g else input_X8_Y13_g when input_X8_Y13_g >= input_X8_Y13_b else input_X8_Y13_b;
output_X8_Y14_gray <= input_X8_Y14_r when input_X8_Y14_r >= input_X8_Y14_b and input_X8_Y14_r >= input_X8_Y14_g else input_X8_Y14_g when input_X8_Y14_g >= input_X8_Y14_b else input_X8_Y14_b;
output_X8_Y15_gray <= input_X8_Y15_r when input_X8_Y15_r >= input_X8_Y15_b and input_X8_Y15_r >= input_X8_Y15_g else input_X8_Y15_g when input_X8_Y15_g >= input_X8_Y15_b else input_X8_Y15_b;
output_X9_Y0_gray <= input_X9_Y0_r when input_X9_Y0_r >= input_X9_Y0_b and input_X9_Y0_r >= input_X9_Y0_g else input_X9_Y0_g when input_X9_Y0_g >= input_X9_Y0_b else input_X9_Y0_b;
output_X9_Y1_gray <= input_X9_Y1_r when input_X9_Y1_r >= input_X9_Y1_b and input_X9_Y1_r >= input_X9_Y1_g else input_X9_Y1_g when input_X9_Y1_g >= input_X9_Y1_b else input_X9_Y1_b;
output_X9_Y2_gray <= input_X9_Y2_r when input_X9_Y2_r >= input_X9_Y2_b and input_X9_Y2_r >= input_X9_Y2_g else input_X9_Y2_g when input_X9_Y2_g >= input_X9_Y2_b else input_X9_Y2_b;
output_X9_Y3_gray <= input_X9_Y3_r when input_X9_Y3_r >= input_X9_Y3_b and input_X9_Y3_r >= input_X9_Y3_g else input_X9_Y3_g when input_X9_Y3_g >= input_X9_Y3_b else input_X9_Y3_b;
output_X9_Y4_gray <= input_X9_Y4_r when input_X9_Y4_r >= input_X9_Y4_b and input_X9_Y4_r >= input_X9_Y4_g else input_X9_Y4_g when input_X9_Y4_g >= input_X9_Y4_b else input_X9_Y4_b;
output_X9_Y5_gray <= input_X9_Y5_r when input_X9_Y5_r >= input_X9_Y5_b and input_X9_Y5_r >= input_X9_Y5_g else input_X9_Y5_g when input_X9_Y5_g >= input_X9_Y5_b else input_X9_Y5_b;
output_X9_Y6_gray <= input_X9_Y6_r when input_X9_Y6_r >= input_X9_Y6_b and input_X9_Y6_r >= input_X9_Y6_g else input_X9_Y6_g when input_X9_Y6_g >= input_X9_Y6_b else input_X9_Y6_b;
output_X9_Y7_gray <= input_X9_Y7_r when input_X9_Y7_r >= input_X9_Y7_b and input_X9_Y7_r >= input_X9_Y7_g else input_X9_Y7_g when input_X9_Y7_g >= input_X9_Y7_b else input_X9_Y7_b;
output_X9_Y8_gray <= input_X9_Y8_r when input_X9_Y8_r >= input_X9_Y8_b and input_X9_Y8_r >= input_X9_Y8_g else input_X9_Y8_g when input_X9_Y8_g >= input_X9_Y8_b else input_X9_Y8_b;
output_X9_Y9_gray <= input_X9_Y9_r when input_X9_Y9_r >= input_X9_Y9_b and input_X9_Y9_r >= input_X9_Y9_g else input_X9_Y9_g when input_X9_Y9_g >= input_X9_Y9_b else input_X9_Y9_b;
output_X9_Y10_gray <= input_X9_Y10_r when input_X9_Y10_r >= input_X9_Y10_b and input_X9_Y10_r >= input_X9_Y10_g else input_X9_Y10_g when input_X9_Y10_g >= input_X9_Y10_b else input_X9_Y10_b;
output_X9_Y11_gray <= input_X9_Y11_r when input_X9_Y11_r >= input_X9_Y11_b and input_X9_Y11_r >= input_X9_Y11_g else input_X9_Y11_g when input_X9_Y11_g >= input_X9_Y11_b else input_X9_Y11_b;
output_X9_Y12_gray <= input_X9_Y12_r when input_X9_Y12_r >= input_X9_Y12_b and input_X9_Y12_r >= input_X9_Y12_g else input_X9_Y12_g when input_X9_Y12_g >= input_X9_Y12_b else input_X9_Y12_b;
output_X9_Y13_gray <= input_X9_Y13_r when input_X9_Y13_r >= input_X9_Y13_b and input_X9_Y13_r >= input_X9_Y13_g else input_X9_Y13_g when input_X9_Y13_g >= input_X9_Y13_b else input_X9_Y13_b;
output_X9_Y14_gray <= input_X9_Y14_r when input_X9_Y14_r >= input_X9_Y14_b and input_X9_Y14_r >= input_X9_Y14_g else input_X9_Y14_g when input_X9_Y14_g >= input_X9_Y14_b else input_X9_Y14_b;
output_X9_Y15_gray <= input_X9_Y15_r when input_X9_Y15_r >= input_X9_Y15_b and input_X9_Y15_r >= input_X9_Y15_g else input_X9_Y15_g when input_X9_Y15_g >= input_X9_Y15_b else input_X9_Y15_b;
output_X10_Y0_gray <= input_X10_Y0_r when input_X10_Y0_r >= input_X10_Y0_b and input_X10_Y0_r >= input_X10_Y0_g else input_X10_Y0_g when input_X10_Y0_g >= input_X10_Y0_b else input_X10_Y0_b;
output_X10_Y1_gray <= input_X10_Y1_r when input_X10_Y1_r >= input_X10_Y1_b and input_X10_Y1_r >= input_X10_Y1_g else input_X10_Y1_g when input_X10_Y1_g >= input_X10_Y1_b else input_X10_Y1_b;
output_X10_Y2_gray <= input_X10_Y2_r when input_X10_Y2_r >= input_X10_Y2_b and input_X10_Y2_r >= input_X10_Y2_g else input_X10_Y2_g when input_X10_Y2_g >= input_X10_Y2_b else input_X10_Y2_b;
output_X10_Y3_gray <= input_X10_Y3_r when input_X10_Y3_r >= input_X10_Y3_b and input_X10_Y3_r >= input_X10_Y3_g else input_X10_Y3_g when input_X10_Y3_g >= input_X10_Y3_b else input_X10_Y3_b;
output_X10_Y4_gray <= input_X10_Y4_r when input_X10_Y4_r >= input_X10_Y4_b and input_X10_Y4_r >= input_X10_Y4_g else input_X10_Y4_g when input_X10_Y4_g >= input_X10_Y4_b else input_X10_Y4_b;
output_X10_Y5_gray <= input_X10_Y5_r when input_X10_Y5_r >= input_X10_Y5_b and input_X10_Y5_r >= input_X10_Y5_g else input_X10_Y5_g when input_X10_Y5_g >= input_X10_Y5_b else input_X10_Y5_b;
output_X10_Y6_gray <= input_X10_Y6_r when input_X10_Y6_r >= input_X10_Y6_b and input_X10_Y6_r >= input_X10_Y6_g else input_X10_Y6_g when input_X10_Y6_g >= input_X10_Y6_b else input_X10_Y6_b;
output_X10_Y7_gray <= input_X10_Y7_r when input_X10_Y7_r >= input_X10_Y7_b and input_X10_Y7_r >= input_X10_Y7_g else input_X10_Y7_g when input_X10_Y7_g >= input_X10_Y7_b else input_X10_Y7_b;
output_X10_Y8_gray <= input_X10_Y8_r when input_X10_Y8_r >= input_X10_Y8_b and input_X10_Y8_r >= input_X10_Y8_g else input_X10_Y8_g when input_X10_Y8_g >= input_X10_Y8_b else input_X10_Y8_b;
output_X10_Y9_gray <= input_X10_Y9_r when input_X10_Y9_r >= input_X10_Y9_b and input_X10_Y9_r >= input_X10_Y9_g else input_X10_Y9_g when input_X10_Y9_g >= input_X10_Y9_b else input_X10_Y9_b;
output_X10_Y10_gray <= input_X10_Y10_r when input_X10_Y10_r >= input_X10_Y10_b and input_X10_Y10_r >= input_X10_Y10_g else input_X10_Y10_g when input_X10_Y10_g >= input_X10_Y10_b else input_X10_Y10_b;
output_X10_Y11_gray <= input_X10_Y11_r when input_X10_Y11_r >= input_X10_Y11_b and input_X10_Y11_r >= input_X10_Y11_g else input_X10_Y11_g when input_X10_Y11_g >= input_X10_Y11_b else input_X10_Y11_b;
output_X10_Y12_gray <= input_X10_Y12_r when input_X10_Y12_r >= input_X10_Y12_b and input_X10_Y12_r >= input_X10_Y12_g else input_X10_Y12_g when input_X10_Y12_g >= input_X10_Y12_b else input_X10_Y12_b;
output_X10_Y13_gray <= input_X10_Y13_r when input_X10_Y13_r >= input_X10_Y13_b and input_X10_Y13_r >= input_X10_Y13_g else input_X10_Y13_g when input_X10_Y13_g >= input_X10_Y13_b else input_X10_Y13_b;
output_X10_Y14_gray <= input_X10_Y14_r when input_X10_Y14_r >= input_X10_Y14_b and input_X10_Y14_r >= input_X10_Y14_g else input_X10_Y14_g when input_X10_Y14_g >= input_X10_Y14_b else input_X10_Y14_b;
output_X10_Y15_gray <= input_X10_Y15_r when input_X10_Y15_r >= input_X10_Y15_b and input_X10_Y15_r >= input_X10_Y15_g else input_X10_Y15_g when input_X10_Y15_g >= input_X10_Y15_b else input_X10_Y15_b;
output_X11_Y0_gray <= input_X11_Y0_r when input_X11_Y0_r >= input_X11_Y0_b and input_X11_Y0_r >= input_X11_Y0_g else input_X11_Y0_g when input_X11_Y0_g >= input_X11_Y0_b else input_X11_Y0_b;
output_X11_Y1_gray <= input_X11_Y1_r when input_X11_Y1_r >= input_X11_Y1_b and input_X11_Y1_r >= input_X11_Y1_g else input_X11_Y1_g when input_X11_Y1_g >= input_X11_Y1_b else input_X11_Y1_b;
output_X11_Y2_gray <= input_X11_Y2_r when input_X11_Y2_r >= input_X11_Y2_b and input_X11_Y2_r >= input_X11_Y2_g else input_X11_Y2_g when input_X11_Y2_g >= input_X11_Y2_b else input_X11_Y2_b;
output_X11_Y3_gray <= input_X11_Y3_r when input_X11_Y3_r >= input_X11_Y3_b and input_X11_Y3_r >= input_X11_Y3_g else input_X11_Y3_g when input_X11_Y3_g >= input_X11_Y3_b else input_X11_Y3_b;
output_X11_Y4_gray <= input_X11_Y4_r when input_X11_Y4_r >= input_X11_Y4_b and input_X11_Y4_r >= input_X11_Y4_g else input_X11_Y4_g when input_X11_Y4_g >= input_X11_Y4_b else input_X11_Y4_b;
output_X11_Y5_gray <= input_X11_Y5_r when input_X11_Y5_r >= input_X11_Y5_b and input_X11_Y5_r >= input_X11_Y5_g else input_X11_Y5_g when input_X11_Y5_g >= input_X11_Y5_b else input_X11_Y5_b;
output_X11_Y6_gray <= input_X11_Y6_r when input_X11_Y6_r >= input_X11_Y6_b and input_X11_Y6_r >= input_X11_Y6_g else input_X11_Y6_g when input_X11_Y6_g >= input_X11_Y6_b else input_X11_Y6_b;
output_X11_Y7_gray <= input_X11_Y7_r when input_X11_Y7_r >= input_X11_Y7_b and input_X11_Y7_r >= input_X11_Y7_g else input_X11_Y7_g when input_X11_Y7_g >= input_X11_Y7_b else input_X11_Y7_b;
output_X11_Y8_gray <= input_X11_Y8_r when input_X11_Y8_r >= input_X11_Y8_b and input_X11_Y8_r >= input_X11_Y8_g else input_X11_Y8_g when input_X11_Y8_g >= input_X11_Y8_b else input_X11_Y8_b;
output_X11_Y9_gray <= input_X11_Y9_r when input_X11_Y9_r >= input_X11_Y9_b and input_X11_Y9_r >= input_X11_Y9_g else input_X11_Y9_g when input_X11_Y9_g >= input_X11_Y9_b else input_X11_Y9_b;
output_X11_Y10_gray <= input_X11_Y10_r when input_X11_Y10_r >= input_X11_Y10_b and input_X11_Y10_r >= input_X11_Y10_g else input_X11_Y10_g when input_X11_Y10_g >= input_X11_Y10_b else input_X11_Y10_b;
output_X11_Y11_gray <= input_X11_Y11_r when input_X11_Y11_r >= input_X11_Y11_b and input_X11_Y11_r >= input_X11_Y11_g else input_X11_Y11_g when input_X11_Y11_g >= input_X11_Y11_b else input_X11_Y11_b;
output_X11_Y12_gray <= input_X11_Y12_r when input_X11_Y12_r >= input_X11_Y12_b and input_X11_Y12_r >= input_X11_Y12_g else input_X11_Y12_g when input_X11_Y12_g >= input_X11_Y12_b else input_X11_Y12_b;
output_X11_Y13_gray <= input_X11_Y13_r when input_X11_Y13_r >= input_X11_Y13_b and input_X11_Y13_r >= input_X11_Y13_g else input_X11_Y13_g when input_X11_Y13_g >= input_X11_Y13_b else input_X11_Y13_b;
output_X11_Y14_gray <= input_X11_Y14_r when input_X11_Y14_r >= input_X11_Y14_b and input_X11_Y14_r >= input_X11_Y14_g else input_X11_Y14_g when input_X11_Y14_g >= input_X11_Y14_b else input_X11_Y14_b;
output_X11_Y15_gray <= input_X11_Y15_r when input_X11_Y15_r >= input_X11_Y15_b and input_X11_Y15_r >= input_X11_Y15_g else input_X11_Y15_g when input_X11_Y15_g >= input_X11_Y15_b else input_X11_Y15_b;
output_X12_Y0_gray <= input_X12_Y0_r when input_X12_Y0_r >= input_X12_Y0_b and input_X12_Y0_r >= input_X12_Y0_g else input_X12_Y0_g when input_X12_Y0_g >= input_X12_Y0_b else input_X12_Y0_b;
output_X12_Y1_gray <= input_X12_Y1_r when input_X12_Y1_r >= input_X12_Y1_b and input_X12_Y1_r >= input_X12_Y1_g else input_X12_Y1_g when input_X12_Y1_g >= input_X12_Y1_b else input_X12_Y1_b;
output_X12_Y2_gray <= input_X12_Y2_r when input_X12_Y2_r >= input_X12_Y2_b and input_X12_Y2_r >= input_X12_Y2_g else input_X12_Y2_g when input_X12_Y2_g >= input_X12_Y2_b else input_X12_Y2_b;
output_X12_Y3_gray <= input_X12_Y3_r when input_X12_Y3_r >= input_X12_Y3_b and input_X12_Y3_r >= input_X12_Y3_g else input_X12_Y3_g when input_X12_Y3_g >= input_X12_Y3_b else input_X12_Y3_b;
output_X12_Y4_gray <= input_X12_Y4_r when input_X12_Y4_r >= input_X12_Y4_b and input_X12_Y4_r >= input_X12_Y4_g else input_X12_Y4_g when input_X12_Y4_g >= input_X12_Y4_b else input_X12_Y4_b;
output_X12_Y5_gray <= input_X12_Y5_r when input_X12_Y5_r >= input_X12_Y5_b and input_X12_Y5_r >= input_X12_Y5_g else input_X12_Y5_g when input_X12_Y5_g >= input_X12_Y5_b else input_X12_Y5_b;
output_X12_Y6_gray <= input_X12_Y6_r when input_X12_Y6_r >= input_X12_Y6_b and input_X12_Y6_r >= input_X12_Y6_g else input_X12_Y6_g when input_X12_Y6_g >= input_X12_Y6_b else input_X12_Y6_b;
output_X12_Y7_gray <= input_X12_Y7_r when input_X12_Y7_r >= input_X12_Y7_b and input_X12_Y7_r >= input_X12_Y7_g else input_X12_Y7_g when input_X12_Y7_g >= input_X12_Y7_b else input_X12_Y7_b;
output_X12_Y8_gray <= input_X12_Y8_r when input_X12_Y8_r >= input_X12_Y8_b and input_X12_Y8_r >= input_X12_Y8_g else input_X12_Y8_g when input_X12_Y8_g >= input_X12_Y8_b else input_X12_Y8_b;
output_X12_Y9_gray <= input_X12_Y9_r when input_X12_Y9_r >= input_X12_Y9_b and input_X12_Y9_r >= input_X12_Y9_g else input_X12_Y9_g when input_X12_Y9_g >= input_X12_Y9_b else input_X12_Y9_b;
output_X12_Y10_gray <= input_X12_Y10_r when input_X12_Y10_r >= input_X12_Y10_b and input_X12_Y10_r >= input_X12_Y10_g else input_X12_Y10_g when input_X12_Y10_g >= input_X12_Y10_b else input_X12_Y10_b;
output_X12_Y11_gray <= input_X12_Y11_r when input_X12_Y11_r >= input_X12_Y11_b and input_X12_Y11_r >= input_X12_Y11_g else input_X12_Y11_g when input_X12_Y11_g >= input_X12_Y11_b else input_X12_Y11_b;
output_X12_Y12_gray <= input_X12_Y12_r when input_X12_Y12_r >= input_X12_Y12_b and input_X12_Y12_r >= input_X12_Y12_g else input_X12_Y12_g when input_X12_Y12_g >= input_X12_Y12_b else input_X12_Y12_b;
output_X12_Y13_gray <= input_X12_Y13_r when input_X12_Y13_r >= input_X12_Y13_b and input_X12_Y13_r >= input_X12_Y13_g else input_X12_Y13_g when input_X12_Y13_g >= input_X12_Y13_b else input_X12_Y13_b;
output_X12_Y14_gray <= input_X12_Y14_r when input_X12_Y14_r >= input_X12_Y14_b and input_X12_Y14_r >= input_X12_Y14_g else input_X12_Y14_g when input_X12_Y14_g >= input_X12_Y14_b else input_X12_Y14_b;
output_X12_Y15_gray <= input_X12_Y15_r when input_X12_Y15_r >= input_X12_Y15_b and input_X12_Y15_r >= input_X12_Y15_g else input_X12_Y15_g when input_X12_Y15_g >= input_X12_Y15_b else input_X12_Y15_b;
output_X13_Y0_gray <= input_X13_Y0_r when input_X13_Y0_r >= input_X13_Y0_b and input_X13_Y0_r >= input_X13_Y0_g else input_X13_Y0_g when input_X13_Y0_g >= input_X13_Y0_b else input_X13_Y0_b;
output_X13_Y1_gray <= input_X13_Y1_r when input_X13_Y1_r >= input_X13_Y1_b and input_X13_Y1_r >= input_X13_Y1_g else input_X13_Y1_g when input_X13_Y1_g >= input_X13_Y1_b else input_X13_Y1_b;
output_X13_Y2_gray <= input_X13_Y2_r when input_X13_Y2_r >= input_X13_Y2_b and input_X13_Y2_r >= input_X13_Y2_g else input_X13_Y2_g when input_X13_Y2_g >= input_X13_Y2_b else input_X13_Y2_b;
output_X13_Y3_gray <= input_X13_Y3_r when input_X13_Y3_r >= input_X13_Y3_b and input_X13_Y3_r >= input_X13_Y3_g else input_X13_Y3_g when input_X13_Y3_g >= input_X13_Y3_b else input_X13_Y3_b;
output_X13_Y4_gray <= input_X13_Y4_r when input_X13_Y4_r >= input_X13_Y4_b and input_X13_Y4_r >= input_X13_Y4_g else input_X13_Y4_g when input_X13_Y4_g >= input_X13_Y4_b else input_X13_Y4_b;
output_X13_Y5_gray <= input_X13_Y5_r when input_X13_Y5_r >= input_X13_Y5_b and input_X13_Y5_r >= input_X13_Y5_g else input_X13_Y5_g when input_X13_Y5_g >= input_X13_Y5_b else input_X13_Y5_b;
output_X13_Y6_gray <= input_X13_Y6_r when input_X13_Y6_r >= input_X13_Y6_b and input_X13_Y6_r >= input_X13_Y6_g else input_X13_Y6_g when input_X13_Y6_g >= input_X13_Y6_b else input_X13_Y6_b;
output_X13_Y7_gray <= input_X13_Y7_r when input_X13_Y7_r >= input_X13_Y7_b and input_X13_Y7_r >= input_X13_Y7_g else input_X13_Y7_g when input_X13_Y7_g >= input_X13_Y7_b else input_X13_Y7_b;
output_X13_Y8_gray <= input_X13_Y8_r when input_X13_Y8_r >= input_X13_Y8_b and input_X13_Y8_r >= input_X13_Y8_g else input_X13_Y8_g when input_X13_Y8_g >= input_X13_Y8_b else input_X13_Y8_b;
output_X13_Y9_gray <= input_X13_Y9_r when input_X13_Y9_r >= input_X13_Y9_b and input_X13_Y9_r >= input_X13_Y9_g else input_X13_Y9_g when input_X13_Y9_g >= input_X13_Y9_b else input_X13_Y9_b;
output_X13_Y10_gray <= input_X13_Y10_r when input_X13_Y10_r >= input_X13_Y10_b and input_X13_Y10_r >= input_X13_Y10_g else input_X13_Y10_g when input_X13_Y10_g >= input_X13_Y10_b else input_X13_Y10_b;
output_X13_Y11_gray <= input_X13_Y11_r when input_X13_Y11_r >= input_X13_Y11_b and input_X13_Y11_r >= input_X13_Y11_g else input_X13_Y11_g when input_X13_Y11_g >= input_X13_Y11_b else input_X13_Y11_b;
output_X13_Y12_gray <= input_X13_Y12_r when input_X13_Y12_r >= input_X13_Y12_b and input_X13_Y12_r >= input_X13_Y12_g else input_X13_Y12_g when input_X13_Y12_g >= input_X13_Y12_b else input_X13_Y12_b;
output_X13_Y13_gray <= input_X13_Y13_r when input_X13_Y13_r >= input_X13_Y13_b and input_X13_Y13_r >= input_X13_Y13_g else input_X13_Y13_g when input_X13_Y13_g >= input_X13_Y13_b else input_X13_Y13_b;
output_X13_Y14_gray <= input_X13_Y14_r when input_X13_Y14_r >= input_X13_Y14_b and input_X13_Y14_r >= input_X13_Y14_g else input_X13_Y14_g when input_X13_Y14_g >= input_X13_Y14_b else input_X13_Y14_b;
output_X13_Y15_gray <= input_X13_Y15_r when input_X13_Y15_r >= input_X13_Y15_b and input_X13_Y15_r >= input_X13_Y15_g else input_X13_Y15_g when input_X13_Y15_g >= input_X13_Y15_b else input_X13_Y15_b;
output_X14_Y0_gray <= input_X14_Y0_r when input_X14_Y0_r >= input_X14_Y0_b and input_X14_Y0_r >= input_X14_Y0_g else input_X14_Y0_g when input_X14_Y0_g >= input_X14_Y0_b else input_X14_Y0_b;
output_X14_Y1_gray <= input_X14_Y1_r when input_X14_Y1_r >= input_X14_Y1_b and input_X14_Y1_r >= input_X14_Y1_g else input_X14_Y1_g when input_X14_Y1_g >= input_X14_Y1_b else input_X14_Y1_b;
output_X14_Y2_gray <= input_X14_Y2_r when input_X14_Y2_r >= input_X14_Y2_b and input_X14_Y2_r >= input_X14_Y2_g else input_X14_Y2_g when input_X14_Y2_g >= input_X14_Y2_b else input_X14_Y2_b;
output_X14_Y3_gray <= input_X14_Y3_r when input_X14_Y3_r >= input_X14_Y3_b and input_X14_Y3_r >= input_X14_Y3_g else input_X14_Y3_g when input_X14_Y3_g >= input_X14_Y3_b else input_X14_Y3_b;
output_X14_Y4_gray <= input_X14_Y4_r when input_X14_Y4_r >= input_X14_Y4_b and input_X14_Y4_r >= input_X14_Y4_g else input_X14_Y4_g when input_X14_Y4_g >= input_X14_Y4_b else input_X14_Y4_b;
output_X14_Y5_gray <= input_X14_Y5_r when input_X14_Y5_r >= input_X14_Y5_b and input_X14_Y5_r >= input_X14_Y5_g else input_X14_Y5_g when input_X14_Y5_g >= input_X14_Y5_b else input_X14_Y5_b;
output_X14_Y6_gray <= input_X14_Y6_r when input_X14_Y6_r >= input_X14_Y6_b and input_X14_Y6_r >= input_X14_Y6_g else input_X14_Y6_g when input_X14_Y6_g >= input_X14_Y6_b else input_X14_Y6_b;
output_X14_Y7_gray <= input_X14_Y7_r when input_X14_Y7_r >= input_X14_Y7_b and input_X14_Y7_r >= input_X14_Y7_g else input_X14_Y7_g when input_X14_Y7_g >= input_X14_Y7_b else input_X14_Y7_b;
output_X14_Y8_gray <= input_X14_Y8_r when input_X14_Y8_r >= input_X14_Y8_b and input_X14_Y8_r >= input_X14_Y8_g else input_X14_Y8_g when input_X14_Y8_g >= input_X14_Y8_b else input_X14_Y8_b;
output_X14_Y9_gray <= input_X14_Y9_r when input_X14_Y9_r >= input_X14_Y9_b and input_X14_Y9_r >= input_X14_Y9_g else input_X14_Y9_g when input_X14_Y9_g >= input_X14_Y9_b else input_X14_Y9_b;
output_X14_Y10_gray <= input_X14_Y10_r when input_X14_Y10_r >= input_X14_Y10_b and input_X14_Y10_r >= input_X14_Y10_g else input_X14_Y10_g when input_X14_Y10_g >= input_X14_Y10_b else input_X14_Y10_b;
output_X14_Y11_gray <= input_X14_Y11_r when input_X14_Y11_r >= input_X14_Y11_b and input_X14_Y11_r >= input_X14_Y11_g else input_X14_Y11_g when input_X14_Y11_g >= input_X14_Y11_b else input_X14_Y11_b;
output_X14_Y12_gray <= input_X14_Y12_r when input_X14_Y12_r >= input_X14_Y12_b and input_X14_Y12_r >= input_X14_Y12_g else input_X14_Y12_g when input_X14_Y12_g >= input_X14_Y12_b else input_X14_Y12_b;
output_X14_Y13_gray <= input_X14_Y13_r when input_X14_Y13_r >= input_X14_Y13_b and input_X14_Y13_r >= input_X14_Y13_g else input_X14_Y13_g when input_X14_Y13_g >= input_X14_Y13_b else input_X14_Y13_b;
output_X14_Y14_gray <= input_X14_Y14_r when input_X14_Y14_r >= input_X14_Y14_b and input_X14_Y14_r >= input_X14_Y14_g else input_X14_Y14_g when input_X14_Y14_g >= input_X14_Y14_b else input_X14_Y14_b;
output_X14_Y15_gray <= input_X14_Y15_r when input_X14_Y15_r >= input_X14_Y15_b and input_X14_Y15_r >= input_X14_Y15_g else input_X14_Y15_g when input_X14_Y15_g >= input_X14_Y15_b else input_X14_Y15_b;
output_X15_Y0_gray <= input_X15_Y0_r when input_X15_Y0_r >= input_X15_Y0_b and input_X15_Y0_r >= input_X15_Y0_g else input_X15_Y0_g when input_X15_Y0_g >= input_X15_Y0_b else input_X15_Y0_b;
output_X15_Y1_gray <= input_X15_Y1_r when input_X15_Y1_r >= input_X15_Y1_b and input_X15_Y1_r >= input_X15_Y1_g else input_X15_Y1_g when input_X15_Y1_g >= input_X15_Y1_b else input_X15_Y1_b;
output_X15_Y2_gray <= input_X15_Y2_r when input_X15_Y2_r >= input_X15_Y2_b and input_X15_Y2_r >= input_X15_Y2_g else input_X15_Y2_g when input_X15_Y2_g >= input_X15_Y2_b else input_X15_Y2_b;
output_X15_Y3_gray <= input_X15_Y3_r when input_X15_Y3_r >= input_X15_Y3_b and input_X15_Y3_r >= input_X15_Y3_g else input_X15_Y3_g when input_X15_Y3_g >= input_X15_Y3_b else input_X15_Y3_b;
output_X15_Y4_gray <= input_X15_Y4_r when input_X15_Y4_r >= input_X15_Y4_b and input_X15_Y4_r >= input_X15_Y4_g else input_X15_Y4_g when input_X15_Y4_g >= input_X15_Y4_b else input_X15_Y4_b;
output_X15_Y5_gray <= input_X15_Y5_r when input_X15_Y5_r >= input_X15_Y5_b and input_X15_Y5_r >= input_X15_Y5_g else input_X15_Y5_g when input_X15_Y5_g >= input_X15_Y5_b else input_X15_Y5_b;
output_X15_Y6_gray <= input_X15_Y6_r when input_X15_Y6_r >= input_X15_Y6_b and input_X15_Y6_r >= input_X15_Y6_g else input_X15_Y6_g when input_X15_Y6_g >= input_X15_Y6_b else input_X15_Y6_b;
output_X15_Y7_gray <= input_X15_Y7_r when input_X15_Y7_r >= input_X15_Y7_b and input_X15_Y7_r >= input_X15_Y7_g else input_X15_Y7_g when input_X15_Y7_g >= input_X15_Y7_b else input_X15_Y7_b;
output_X15_Y8_gray <= input_X15_Y8_r when input_X15_Y8_r >= input_X15_Y8_b and input_X15_Y8_r >= input_X15_Y8_g else input_X15_Y8_g when input_X15_Y8_g >= input_X15_Y8_b else input_X15_Y8_b;
output_X15_Y9_gray <= input_X15_Y9_r when input_X15_Y9_r >= input_X15_Y9_b and input_X15_Y9_r >= input_X15_Y9_g else input_X15_Y9_g when input_X15_Y9_g >= input_X15_Y9_b else input_X15_Y9_b;
output_X15_Y10_gray <= input_X15_Y10_r when input_X15_Y10_r >= input_X15_Y10_b and input_X15_Y10_r >= input_X15_Y10_g else input_X15_Y10_g when input_X15_Y10_g >= input_X15_Y10_b else input_X15_Y10_b;
output_X15_Y11_gray <= input_X15_Y11_r when input_X15_Y11_r >= input_X15_Y11_b and input_X15_Y11_r >= input_X15_Y11_g else input_X15_Y11_g when input_X15_Y11_g >= input_X15_Y11_b else input_X15_Y11_b;
output_X15_Y12_gray <= input_X15_Y12_r when input_X15_Y12_r >= input_X15_Y12_b and input_X15_Y12_r >= input_X15_Y12_g else input_X15_Y12_g when input_X15_Y12_g >= input_X15_Y12_b else input_X15_Y12_b;
output_X15_Y13_gray <= input_X15_Y13_r when input_X15_Y13_r >= input_X15_Y13_b and input_X15_Y13_r >= input_X15_Y13_g else input_X15_Y13_g when input_X15_Y13_g >= input_X15_Y13_b else input_X15_Y13_b;
output_X15_Y14_gray <= input_X15_Y14_r when input_X15_Y14_r >= input_X15_Y14_b and input_X15_Y14_r >= input_X15_Y14_g else input_X15_Y14_g when input_X15_Y14_g >= input_X15_Y14_b else input_X15_Y14_b;
output_X15_Y15_gray <= input_X15_Y15_r when input_X15_Y15_r >= input_X15_Y15_b and input_X15_Y15_r >= input_X15_Y15_g else input_X15_Y15_g when input_X15_Y15_g >= input_X15_Y15_b else input_X15_Y15_b;


end Behavioral;


